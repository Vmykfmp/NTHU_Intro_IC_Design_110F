* SPICE NETLIST
***************************************
*HW2_Inverter_Chain_postsim
.lib 'cic018.l' TT
.temp 25
.unprot
.inc "IC.pex.spi"
.option post

*Voltage
V1 VDD 0 1.8
V2 GND 0 0
VVIN_pulse Vin GND pulse 0 1.8 10n 1n 1n 4n 10n

*Capacitor
CL Vout GND 10pF

*Circuit
x1 Vin GND VDD Vout IC

*simulation setup
.Tran 1ps 50ns
.MEAS tran TpHL_Vout trig V(Vin) val=0.9 td=0 rise=1 targ V(Vout) val=0.9 fall=1
.MEAS tran TpLH_Vout trig V(Vin) val=0.9 td=0 fall=1 targ V(Vout) val=0.9 rise=1

.SUBCKT L POS NEG
.ENDS
.end
***************************************
.SUBCKT IC Vin GND VDD Vout
** N=6 EP=4 IP=0 FDC=94
M0 2 Vin GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=4765 $Y=-166 $D=0
M1 3 2 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=6325 $Y=-166 $D=0
M2 GND 2 3 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=7015 $Y=-166 $D=0
M3 3 2 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=7705 $Y=-166 $D=0
M4 GND 2 3 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=8395 $Y=-166 $D=0
M5 3 2 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=9085 $Y=-166 $D=0
M6 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=10645 $Y=-166 $D=0
M7 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=11335 $Y=-166 $D=0
M8 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=12025 $Y=-166 $D=0
M9 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=12715 $Y=-166 $D=0
M10 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=13405 $Y=-166 $D=0
M11 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=14095 $Y=-166 $D=0
M12 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=14785 $Y=-166 $D=0
M13 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=15475 $Y=-166 $D=0
M14 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=16165 $Y=-166 $D=0
M15 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=16855 $Y=-166 $D=0
M16 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=17545 $Y=-166 $D=0
M17 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=18235 $Y=-166 $D=0
M18 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=18925 $Y=-166 $D=0
M19 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=19615 $Y=-166 $D=0
M20 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=20305 $Y=-166 $D=0
M21 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=20995 $Y=-166 $D=0
M22 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=21685 $Y=-166 $D=0
M23 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=22375 $Y=-166 $D=0
M24 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=23065 $Y=-166 $D=0
M25 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=23755 $Y=-166 $D=0
M26 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=24445 $Y=-166 $D=0
M27 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=25135 $Y=-166 $D=0
M28 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=25825 $Y=-166 $D=0
M29 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=26515 $Y=-166 $D=0
M30 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=27205 $Y=-166 $D=0
M31 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=27895 $Y=-166 $D=0
M32 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=28585 $Y=-166 $D=0
M33 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=29275 $Y=-166 $D=0
M34 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=29965 $Y=-166 $D=0
M35 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=30655 $Y=-166 $D=0
M36 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=31345 $Y=-166 $D=0
M37 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=32035 $Y=-166 $D=0
M38 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=32725 $Y=-166 $D=0
M39 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=33415 $Y=-166 $D=0
M40 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=34105 $Y=-166 $D=0
M41 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=34795 $Y=-166 $D=0
M42 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=35485 $Y=-166 $D=0
M43 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=36175 $Y=-166 $D=0
M44 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=36865 $Y=-166 $D=0
M45 GND 3 Vout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=37555 $Y=-166 $D=0
M46 Vout 3 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=38245 $Y=-166 $D=0
M47 2 Vin VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=9.0454e-13 PD=2.826e-06 PS=2.826e-06 $X=4765 $Y=1334 $D=1
M48 3 2 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=6325 $Y=1334 $D=1
M49 VDD 2 3 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=7015 $Y=1334 $D=1
M50 3 2 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=7705 $Y=1334 $D=1
M51 VDD 2 3 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=8395 $Y=1334 $D=1
M52 3 2 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=9085 $Y=1334 $D=1
M53 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=10645 $Y=1334 $D=1
M54 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=11335 $Y=1334 $D=1
M55 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=12025 $Y=1334 $D=1
M56 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=12715 $Y=1334 $D=1
M57 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=13405 $Y=1334 $D=1
M58 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=14095 $Y=1334 $D=1
M59 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=14785 $Y=1334 $D=1
M60 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=15475 $Y=1334 $D=1
M61 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=16165 $Y=1334 $D=1
M62 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=16855 $Y=1334 $D=1
M63 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=17545 $Y=1334 $D=1
M64 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=18235 $Y=1334 $D=1
M65 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=18925 $Y=1334 $D=1
M66 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=19615 $Y=1334 $D=1
M67 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=20305 $Y=1334 $D=1
M68 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=20995 $Y=1334 $D=1
M69 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=21685 $Y=1334 $D=1
M70 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=22375 $Y=1334 $D=1
M71 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=23065 $Y=1334 $D=1
M72 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=23755 $Y=1334 $D=1
M73 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=24445 $Y=1334 $D=1
M74 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=25135 $Y=1334 $D=1
M75 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=25825 $Y=1334 $D=1
M76 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=26515 $Y=1334 $D=1
M77 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=27205 $Y=1334 $D=1
M78 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=27895 $Y=1334 $D=1
M79 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=28585 $Y=1334 $D=1
M80 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=29275 $Y=1334 $D=1
M81 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=29965 $Y=1334 $D=1
M82 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=30655 $Y=1334 $D=1
M83 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=31345 $Y=1334 $D=1
M84 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=32035 $Y=1334 $D=1
M85 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=32725 $Y=1334 $D=1
M86 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=33415 $Y=1334 $D=1
M87 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=34105 $Y=1334 $D=1
M88 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=34795 $Y=1334 $D=1
M89 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=35485 $Y=1334 $D=1
M90 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=36175 $Y=1334 $D=1
M91 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=36865 $Y=1334 $D=1
M92 VDD 3 Vout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=37555 $Y=1334 $D=1
M93 Vout 3 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=38245 $Y=1334 $D=1
.ENDS
***************************************
