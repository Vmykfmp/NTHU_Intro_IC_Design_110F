* File: top.pex.spi
* Created: Tue Jan 18 17:29:49 2022
* Program "Calibre xRC"
* Version "v2021.1_33.19"
* 
.include "top.pex.spi.pex"
.subckt top  CLK VREF VDD VSS DOUT<0> DOUT<1> A<2> A<5> A<6> A<7> A<8> A<1> A<0>
+ A<3> A<4>
* 
* A<4>	A<4>
* A<3>	A<3>
* A<0>	A<0>
* A<1>	A<1>
* A<8>	A<8>
* A<7>	A<7>
* A<6>	A<6>
* A<5>	A<5>
* A<2>	A<2>
* DOUT<1>	DOUT<1>
* DOUT<0>	DOUT<0>
* VSS	VSS
* VDD	VDD
* VREF	VREF
* CLK	CLK
mXDFF_Timing_control/XI9/XI2/MM5
+ N_XDFF_TIMING_CONTROL/XI9/XI2/NET41_XDFF_Timing_control/XI9/XI2/MM5_d
+ N_CLK_XDFF_Timing_control/XI9/XI2/MM5_g
+ N_VSS_XDFF_Timing_control/XI9/XI2/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b
+ N_18 L=6e-07 W=5e-07 AD=2.95e-13 AS=2.45e-13 PD=1.68e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI2/MM6
+ N_XDFF_TIMING_CONTROL/XI9/XI2/NET37_XDFF_Timing_control/XI9/XI2/MM6_d
+ N_XDFF_TIMING_CONTROL/XI9/XI2/NET41_XDFF_Timing_control/XI9/XI2/MM6_g
+ N_VSS_XDFF_Timing_control/XI9/XI2/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b
+ N_18 L=6e-07 W=5e-07 AD=2.95e-13 AS=2.45e-13 PD=1.68e-06 PS=1.48e-06
mXYDec/XI17/MN N_XYDEC/NET22_XYDec/XI17/MN_d N_Y_SEL_FF<0>_XYDec/XI17/MN_g
+ N_VSS_XYDec/XI17/MN_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI2/MM7
+ N_XDFF_TIMING_CONTROL/XI9/XI2/NET33_XDFF_Timing_control/XI9/XI2/MM7_d
+ N_XDFF_TIMING_CONTROL/XI9/XI2/NET37_XDFF_Timing_control/XI9/XI2/MM7_g
+ N_VSS_XDFF_Timing_control/XI9/XI2/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b
+ N_18 L=6e-07 W=5e-07 AD=2.95e-13 AS=2.45e-13 PD=1.68e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI2/MM8
+ N_XDFF_TIMING_CONTROL/XI9/NET10_XDFF_Timing_control/XI9/XI2/MM8_d
+ N_XDFF_TIMING_CONTROL/XI9/XI2/NET33_XDFF_Timing_control/XI9/XI2/MM8_g
+ N_VSS_XDFF_Timing_control/XI9/XI2/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b
+ N_18 L=6e-07 W=5e-07 AD=2.95e-13 AS=2.45e-13 PD=1.68e-06 PS=1.48e-06
mXYDec/XI18/MN N_XYDEC/NET18_XYDec/XI18/MN_d N_Y_SEL_FF<1>_XYDec/XI18/MN_g
+ N_VSS_XYDec/XI18/MN_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/MMMa
+ N_XDFF_TIMING_CONTROL/XI9/NET023_XDFF_Timing_control/XI9/MMMa_d
+ N_XDFF_TIMING_CONTROL/XI9/NET10_XDFF_Timing_control/XI9/MMMa_g
+ N_VSS_XDFF_Timing_control/XI9/MMMa_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1e-06 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXYDec/XI19/MN N_XYDEC/NET14_XYDec/XI19/MN_d N_Y_SEL_FF<2>_XYDec/XI19/MN_g
+ N_VSS_XYDec/XI19/MN_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/MMMc
+ N_XDFF_TIMING_CONTROL/XI9/NET013_XDFF_Timing_control/XI9/MMMc_d
+ N_XDFF_TIMING_CONTROL/XI9/NET023_XDFF_Timing_control/XI9/MMMc_g
+ N_VSS_XDFF_Timing_control/XI9/MMMc_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1e-06 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI1/XI2/MM5
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI2/NET41_XDFF_Timing_control/XI9/XI1/XI2/MM5_d
+ N_XDFF_TIMING_CONTROL/XI9/NET013_XDFF_Timing_control/XI9/XI1/XI2/MM5_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI2/MM5_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=6e-07 W=5e-07 AD=2.95e-13
+ AS=2.45e-13 PD=1.68e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI2/MM5
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI2/NET41_XDFF_Timing_control/XI9/XI0/XI2/MM5_d
+ N_CLK_XDFF_Timing_control/XI9/XI0/XI2/MM5_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI2/MM5_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=6e-07 W=5e-07 AD=2.95e-13
+ AS=2.45e-13 PD=1.68e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI1/XI2/MM6
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI2/NET37_XDFF_Timing_control/XI9/XI1/XI2/MM6_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI2/NET41_XDFF_Timing_control/XI9/XI1/XI2/MM6_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI2/MM6_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=6e-07 W=5e-07 AD=2.95e-13
+ AS=2.45e-13 PD=1.68e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI2/MM6
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI2/NET37_XDFF_Timing_control/XI9/XI0/XI2/MM6_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI2/NET41_XDFF_Timing_control/XI9/XI0/XI2/MM6_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI2/MM6_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=6e-07 W=5e-07 AD=2.95e-13
+ AS=2.45e-13 PD=1.68e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI1/XI2/MM7
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI2/NET33_XDFF_Timing_control/XI9/XI1/XI2/MM7_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI2/NET37_XDFF_Timing_control/XI9/XI1/XI2/MM7_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI2/MM7_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=6e-07 W=5e-07 AD=2.95e-13
+ AS=2.45e-13 PD=1.68e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI2/MM7
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI2/NET33_XDFF_Timing_control/XI9/XI0/XI2/MM7_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI2/NET37_XDFF_Timing_control/XI9/XI0/XI2/MM7_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI2/MM7_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=6e-07 W=5e-07 AD=2.95e-13
+ AS=2.45e-13 PD=1.68e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI1/XI2/MM8
+ N_XDFF_TIMING_CONTROL/XI9/XI1/NET011_XDFF_Timing_control/XI9/XI1/XI2/MM8_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI2/NET33_XDFF_Timing_control/XI9/XI1/XI2/MM8_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI2/MM8_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=6e-07 W=5e-07 AD=3e-13 AS=2.45e-13
+ PD=1.7e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI2/MM8
+ N_XDFF_TIMING_CONTROL/XI9/XI0/NET011_XDFF_Timing_control/XI9/XI0/XI2/MM8_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI2/NET33_XDFF_Timing_control/XI9/XI0/XI2/MM8_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI2/MM8_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=6e-07 W=5e-07 AD=3e-13 AS=2.45e-13
+ PD=1.7e-06 PS=1.48e-06
mXYDec/XI21/MM3 N_XYDEC/XI21/NET24_XYDec/XI21/MM3_d N_VDD_XYDec/XI21/MM3_g
+ N_VSS_XYDec/XI21/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXYDec/XI22/MM3 N_XYDEC/XI22/NET24_XYDec/XI22/MM3_d N_VDD_XYDec/XI22/MM3_g
+ N_VSS_XYDec/XI22/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXYDec/XI25/MM3 N_XYDEC/XI25/NET24_XYDec/XI25/MM3_d N_VDD_XYDec/XI25/MM3_g
+ N_VSS_XYDec/XI25/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXYDec/XI26/MM3 N_XYDEC/XI26/NET24_XYDec/XI26/MM3_d N_VDD_XYDec/XI26/MM3_g
+ N_VSS_XYDec/XI26/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXYDec/XI21/MM2 N_XYDEC/XI21/NET28_XYDec/XI21/MM2_d
+ N_Y_SEL_FF<2>_XYDec/XI21/MM2_g N_XYDEC/XI21/NET24_XYDec/XI21/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI22/MM2 N_XYDEC/XI22/NET28_XYDec/XI22/MM2_d
+ N_Y_SEL_FF<2>_XYDec/XI22/MM2_g N_XYDEC/XI22/NET24_XYDec/XI22/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI25/MM2 N_XYDEC/XI25/NET28_XYDec/XI25/MM2_d
+ N_XYDEC/NET14_XYDec/XI25/MM2_g N_XYDEC/XI25/NET24_XYDec/XI25/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI26/MM2 N_XYDEC/XI26/NET28_XYDec/XI26/MM2_d
+ N_XYDEC/NET14_XYDec/XI26/MM2_g N_XYDEC/XI26/NET24_XYDec/XI26/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXDFF_Timing_control/XI9/XI1/XI1/MM5
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET39_XDFF_Timing_control/XI9/XI1/XI1/MM5_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/NET011_XDFF_Timing_control/XI9/XI1/XI1/MM5_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI1/MM5_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI1/MM5
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET39_XDFF_Timing_control/XI9/XI0/XI1/MM5_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/NET011_XDFF_Timing_control/XI9/XI0/XI1/MM5_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI1/MM5_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXYDec/XI21/MM1 N_XYDEC/XI21/NET32_XYDec/XI21/MM1_d
+ N_Y_SEL_FF<1>_XYDec/XI21/MM1_g N_XYDEC/XI21/NET28_XYDec/XI21/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI22/MM1 N_XYDEC/XI22/NET32_XYDec/XI22/MM1_d
+ N_XYDEC/NET18_XYDec/XI22/MM1_g N_XYDEC/XI22/NET28_XYDec/XI22/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI25/MM1 N_XYDEC/XI25/NET32_XYDec/XI25/MM1_d
+ N_Y_SEL_FF<1>_XYDec/XI25/MM1_g N_XYDEC/XI25/NET28_XYDec/XI25/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI26/MM1 N_XYDEC/XI26/NET32_XYDec/XI26/MM1_d
+ N_XYDEC/NET18_XYDec/XI26/MM1_g N_XYDEC/XI26/NET28_XYDec/XI26/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI21/MM0 N_Y_SEL<6>_XYDec/XI21/MM0_d N_XYDEC/NET22_XYDec/XI21/MM0_g
+ N_XYDEC/XI21/NET32_XYDec/XI21/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI22/MM0 N_Y_SEL<5>_XYDec/XI22/MM0_d N_Y_SEL_FF<0>_XYDec/XI22/MM0_g
+ N_XYDEC/XI22/NET32_XYDec/XI22/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI25/MM0 N_Y_SEL<2>_XYDec/XI25/MM0_d N_XYDEC/NET22_XYDec/XI25/MM0_g
+ N_XYDEC/XI25/NET32_XYDec/XI25/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI26/MM0 N_Y_SEL<1>_XYDec/XI26/MM0_d N_Y_SEL_FF<0>_XYDec/XI26/MM0_g
+ N_XYDEC/XI26/NET32_XYDec/XI26/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI20/MM3 N_XYDEC/XI20/NET24_XYDec/XI20/MM3_d N_VDD_XYDec/XI20/MM3_g
+ N_VSS_XYDec/XI20/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXYDec/XI23/MM3 N_XYDEC/XI23/NET24_XYDec/XI23/MM3_d N_VDD_XYDec/XI23/MM3_g
+ N_VSS_XYDec/XI23/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXYDec/XI24/MM3 N_XYDEC/XI24/NET24_XYDec/XI24/MM3_d N_VDD_XYDec/XI24/MM3_g
+ N_VSS_XYDec/XI24/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXYDec/XI27/MM3 N_XYDEC/XI27/NET24_XYDec/XI27/MM3_d N_VDD_XYDec/XI27/MM3_g
+ N_VSS_XYDec/XI27/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI9/XI1/XI1/MM6
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET15_XDFF_Timing_control/XI9/XI1/XI1/MM6_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET39_XDFF_Timing_control/XI9/XI1/XI1/MM6_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI1/MM6_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI1/MM6
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET15_XDFF_Timing_control/XI9/XI0/XI1/MM6_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET39_XDFF_Timing_control/XI9/XI0/XI1/MM6_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI1/MM6_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXYDec/XI20/MM2 N_XYDEC/XI20/NET28_XYDec/XI20/MM2_d
+ N_Y_SEL_FF<2>_XYDec/XI20/MM2_g N_XYDEC/XI20/NET24_XYDec/XI20/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI23/MM2 N_XYDEC/XI23/NET28_XYDec/XI23/MM2_d
+ N_Y_SEL_FF<2>_XYDec/XI23/MM2_g N_XYDEC/XI23/NET24_XYDec/XI23/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI24/MM2 N_XYDEC/XI24/NET28_XYDec/XI24/MM2_d
+ N_XYDEC/NET14_XYDec/XI24/MM2_g N_XYDEC/XI24/NET24_XYDec/XI24/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI27/MM2 N_XYDEC/XI27/NET28_XYDec/XI27/MM2_d
+ N_XYDEC/NET14_XYDec/XI27/MM2_g N_XYDEC/XI27/NET24_XYDec/XI27/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI20/MM1 N_XYDEC/XI20/NET32_XYDec/XI20/MM1_d
+ N_Y_SEL_FF<1>_XYDec/XI20/MM1_g N_XYDEC/XI20/NET28_XYDec/XI20/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI23/MM1 N_XYDEC/XI23/NET32_XYDec/XI23/MM1_d
+ N_XYDEC/NET18_XYDec/XI23/MM1_g N_XYDEC/XI23/NET28_XYDec/XI23/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI24/MM1 N_XYDEC/XI24/NET32_XYDec/XI24/MM1_d
+ N_Y_SEL_FF<1>_XYDec/XI24/MM1_g N_XYDEC/XI24/NET28_XYDec/XI24/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI27/MM1 N_XYDEC/XI27/NET32_XYDec/XI27/MM1_d
+ N_XYDEC/NET18_XYDec/XI27/MM1_g N_XYDEC/XI27/NET28_XYDec/XI27/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI20/MM0 N_Y_SEL<7>_XYDec/XI20/MM0_d N_Y_SEL_FF<0>_XYDec/XI20/MM0_g
+ N_XYDEC/XI20/NET32_XYDec/XI20/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI23/MM0 N_Y_SEL<4>_XYDec/XI23/MM0_d N_XYDEC/NET22_XYDec/XI23/MM0_g
+ N_XYDEC/XI23/NET32_XYDec/XI23/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI24/MM0 N_Y_SEL<3>_XYDec/XI24/MM0_d N_Y_SEL_FF<0>_XYDec/XI24/MM0_g
+ N_XYDEC/XI24/NET32_XYDec/XI24/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI27/MM0 N_Y_SEL<0>_XYDec/XI27/MM0_d N_XYDEC/NET22_XYDec/XI27/MM0_g
+ N_XYDEC/XI27/NET32_XYDec/XI27/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI9/XI1/XI1/MM7
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET31_XDFF_Timing_control/XI9/XI1/XI1/MM7_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET15_XDFF_Timing_control/XI9/XI1/XI1/MM7_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI1/MM7_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI1/MM7
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET31_XDFF_Timing_control/XI9/XI0/XI1/MM7_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET15_XDFF_Timing_control/XI9/XI0/XI1/MM7_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI1/MM7_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI1/XI1/MM8
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET27_XDFF_Timing_control/XI9/XI1/XI1/MM8_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET31_XDFF_Timing_control/XI9/XI1/XI1/MM8_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI1/MM8_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI1/MM8
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET27_XDFF_Timing_control/XI9/XI0/XI1/MM8_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET31_XDFF_Timing_control/XI9/XI0/XI1/MM8_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI1/MM8_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/MM1 N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/MM1_d
+ N_CLK_XDFF_Timing_control/MM1_g N_VSS_XDFF_Timing_control/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI1/XI1/MM9
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET046_XDFF_Timing_control/XI9/XI1/XI1/MM9_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET27_XDFF_Timing_control/XI9/XI1/XI1/MM9_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI1/MM9_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI1/MM9
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET046_XDFF_Timing_control/XI9/XI0/XI1/MM9_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET27_XDFF_Timing_control/XI9/XI0/XI1/MM9_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI1/MM9_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI1/XI1/MMa
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET038_XDFF_Timing_control/XI9/XI1/XI1/MMa_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET046_XDFF_Timing_control/XI9/XI1/XI1/MMa_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI1/MMa_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI1/MMa
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET038_XDFF_Timing_control/XI9/XI0/XI1/MMa_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET046_XDFF_Timing_control/XI9/XI0/XI1/MMa_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI1/MMa_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI1/XI1/MMc
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET034_XDFF_Timing_control/XI9/XI1/XI1/MMc_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET038_XDFF_Timing_control/XI9/XI1/XI1/MMc_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI1/MMc_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI1/MMc
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET034_XDFF_Timing_control/XI9/XI0/XI1/MMc_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET038_XDFF_Timing_control/XI9/XI0/XI1/MMc_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI1/MMc_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI1/XI1/MMe
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET030_XDFF_Timing_control/XI9/XI1/XI1/MMe_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET034_XDFF_Timing_control/XI9/XI1/XI1/MMe_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI1/MMe_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI1/MMe
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET030_XDFF_Timing_control/XI9/XI0/XI1/MMe_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET034_XDFF_Timing_control/XI9/XI0/XI1/MMe_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI1/MMe_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI1/XI1/MMg
+ N_XDFF_TIMING_CONTROL/XI9/XI1/NET6_XDFF_Timing_control/XI9/XI1/XI1/MMg_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET030_XDFF_Timing_control/XI9/XI1/XI1/MMg_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI1/MMg_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI1/MMg
+ N_XDFF_TIMING_CONTROL/XI9/XI0/NET6_XDFF_Timing_control/XI9/XI0/XI1/MMg_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET030_XDFF_Timing_control/XI9/XI0/XI1/MMg_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI1/MMg_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1e-06 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI1/XI0/MM2
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI0/NET10_XDFF_Timing_control/XI9/XI1/XI0/MM2_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/NET011_XDFF_Timing_control/XI9/XI1/XI0/MM2_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI0/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5.2e-07 AD=1.326e-13
+ AS=2.548e-13 PD=5.1e-07 PS=1.5e-06
mXDFF_Timing_control/XI9/XI0/XI0/MM2
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI0/NET10_XDFF_Timing_control/XI9/XI0/XI0/MM2_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/NET011_XDFF_Timing_control/XI9/XI0/XI0/MM2_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI0/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5.2e-07 AD=1.326e-13
+ AS=2.548e-13 PD=5.1e-07 PS=1.5e-06
mXDFF_Timing_control/XI9/XI1/XI0/MM3
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI0/NET055_XDFF_Timing_control/XI9/XI1/XI0/MM3_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/NET6_XDFF_Timing_control/XI9/XI1/XI0/MM3_g
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI0/NET10_XDFF_Timing_control/XI9/XI1/XI0/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5.2e-07 AD=2.548e-13
+ AS=1.326e-13 PD=1.5e-06 PS=5.1e-07
mXDFF_Timing_control/XI9/XI0/XI0/MM3
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI0/NET055_XDFF_Timing_control/XI9/XI0/XI0/MM3_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/NET6_XDFF_Timing_control/XI9/XI0/XI0/MM3_g
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI0/NET10_XDFF_Timing_control/XI9/XI0/XI0/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5.2e-07 AD=2.548e-13
+ AS=1.326e-13 PD=1.5e-06 PS=5.1e-07
mXDFF_Timing_control/XI9/XI1/XI0/MM4
+ N_SAEN_XDFF_Timing_control/XI9/XI1/XI0/MM4_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI0/NET055_XDFF_Timing_control/XI9/XI1/XI0/MM4_g
+ N_VSS_XDFF_Timing_control/XI9/XI1/XI0/MM4_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI0/XI0/MM4
+ N_WL_EN_XDFF_Timing_control/XI9/XI0/XI0/MM4_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI0/NET055_XDFF_Timing_control/XI9/XI0/XI0/MM4_g
+ N_VSS_XDFF_Timing_control/XI9/XI0/XI0/MM4_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI63/MM1 N_XMUX/NET44_XMUX/XI63/MM1_d N_Y_SEL<7>_XMUX/XI63/MM1_g
+ N_VSS_XMUX/XI63/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI62/MM1 N_XMUX/NET068_XMUX/XI62/MM1_d N_Y_SEL<6>_XMUX/XI62/MM1_g
+ N_VSS_XMUX/XI62/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI61/MM1 N_XMUX/NET106_XMUX/XI61/MM1_d N_Y_SEL<5>_XMUX/XI61/MM1_g
+ N_VSS_XMUX/XI61/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI60/MM1 N_XMUX/NET56_XMUX/XI60/MM1_d N_Y_SEL<4>_XMUX/XI60/MM1_g
+ N_VSS_XMUX/XI60/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI59/MM1 N_XMUX/NET154_XMUX/XI59/MM1_d N_Y_SEL<3>_XMUX/XI59/MM1_g
+ N_VSS_XMUX/XI59/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI58/MM1 N_XMUX/NET130_XMUX/XI58/MM1_d N_Y_SEL<2>_XMUX/XI58/MM1_g
+ N_VSS_XMUX/XI58/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI57/MM1 N_XMUX/NET100_XMUX/XI57/MM1_d N_Y_SEL<1>_XMUX/XI57/MM1_g
+ N_VSS_XMUX/XI57/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI56/MM1 N_XMUX/NET044_XMUX/XI56/MM1_d N_Y_SEL<0>_XMUX/XI56/MM1_g
+ N_VSS_XMUX/XI56/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSRL/MM23 N_XSRL/CLKB_XSRL/MM23_d N_SAEN_XSRL/MM23_g N_VSS_XSRL/MM23_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13
+ AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXSA/MM15 N_XSA/NET060_XSA/MM15_d N_DL<0>_XSA/MM15_g N_XSA/NET0108_XSA/MM15_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.28e-13
+ AS=2.45e-13 PD=5.12e-07 PS=1.48e-06
mXSA/MM11 N_O0_XSA/MM11_d N_DOUT_SA<0>_XSA/MM11_g N_XSA/NET060_XSA/MM11_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.28e-13 PD=1.48e-06 PS=5.12e-07
mXMUX/XI40/MM0 N_BL<0>_XMUX/XI40/MM0_d N_XMUX/NET044_XMUX/XI40/MM0_g
+ N_DL<0>_XMUX/XI40/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI41/MM0 N_BL<1>_XMUX/XI41/MM0_d N_XMUX/NET100_XMUX/XI41/MM0_g
+ N_DL<0>_XMUX/XI41/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI42/MM0 N_BL<2>_XMUX/XI42/MM0_d N_XMUX/NET130_XMUX/XI42/MM0_g
+ N_DL<0>_XMUX/XI42/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSA/MM19 N_XSA/NET0108_XSA/MM19_d N_SAEN_XSA/MM19_g N_VSS_XSA/MM19_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXMUX/XI43/MM0 N_BL<3>_XMUX/XI43/MM0_d N_XMUX/NET154_XMUX/XI43/MM0_g
+ N_DL<0>_XMUX/XI43/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI44/MM0 N_BL<4>_XMUX/XI44/MM0_d N_XMUX/NET56_XMUX/XI44/MM0_g
+ N_DL<0>_XMUX/XI44/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI45/MM0 N_BL<5>_XMUX/XI45/MM0_d N_XMUX/NET106_XMUX/XI45/MM0_g
+ N_DL<0>_XMUX/XI45/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSRL/MM20 N_QB<0>_XSRL/MM20_d N_DOUT<0>_XSRL/MM20_g N_VSS_XSRL/MM20_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13
+ AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXSRL/MM44 N_DOUT<0>_XSRL/MM44_d N_XSRL/CLKB_XSRL/MM44_g
+ N_XSRL/NET0180_XSRL/MM44_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=9.5e-07 AD=2.4225e-13 AS=4.655e-13 PD=5.1e-07 PS=1.93e-06
mXSRL/MM21 N_XSRL/SA0_XSRL/MM21_d N_SAEN_XSRL/MM21_g N_DOUT<0>_XSRL/MM21_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13
+ AS=2.4225e-13 PD=1.93e-06 PS=5.1e-07
mXSRL/MM24 N_XSRL/SA0_XSRL/MM24_d N_XSRL/NET088_XSRL/MM24_g N_VSS_XSRL/MM24_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13
+ AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXSRL/MM25 N_XSRL/NET088_XSRL/MM25_d N_DOUT_SA<0>_XSRL/MM25_g N_VSS_XSRL/MM25_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13
+ AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXMUX/XI46/MM0 N_BL<6>_XMUX/XI46/MM0_d N_XMUX/NET068_XMUX/XI46/MM0_g
+ N_DL<0>_XMUX/XI46/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSA/MM16 N_XSA/NET087_XSA/MM16_d N_VREF_XSA/MM16_g N_XSA/NET0108_XSA/MM16_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.28e-13
+ AS=2.45e-13 PD=5.12e-07 PS=1.48e-06
mXSA/MM13 N_DOUT_SA<0>_XSA/MM13_d N_O0_XSA/MM13_g N_XSA/NET087_XSA/MM13_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.28e-13 PD=1.48e-06 PS=5.12e-07
mXSRL/MM19 N_XSRL/NET0180_XSRL/MM19_d N_QB<0>_XSRL/MM19_g N_VSS_XSRL/MM19_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXMUX/XI47/MM0 N_BL<7>_XMUX/XI47/MM0_d N_XMUX/NET44_XMUX/XI47/MM0_g
+ N_DL<0>_XMUX/XI47/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSA/MM5 N_XSA/NET09_XSA/MM5_d N_DL<1>_XSA/MM5_g N_XSA/NET012_XSA/MM5_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.28e-13
+ AS=2.45e-13 PD=5.12e-07 PS=1.48e-06
mXSA/MM1 N_O1_XSA/MM1_d N_DOUT_SA<1>_XSA/MM1_g N_XSA/NET09_XSA/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.28e-13 PD=1.48e-06 PS=5.12e-07
mXMUX/XI55/MM0 N_BL<8>_XMUX/XI55/MM0_d N_XMUX/NET044_XMUX/XI55/MM0_g
+ N_DL<1>_XMUX/XI55/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSRL/MM56 N_QB<1>_XSRL/MM56_d N_DOUT<1>_XSRL/MM56_g N_VSS_XSRL/MM56_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13
+ AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXSRL/MM55 N_XSRL/NET0178_XSRL/MM55_d N_QB<1>_XSRL/MM55_g N_VSS_XSRL/MM55_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXSRL/MM54 N_DOUT<1>_XSRL/MM54_d N_XSRL/CLKB_XSRL/MM54_g
+ N_XSRL/NET0178_XSRL/MM54_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=9.5e-07 AD=2.4225e-13 AS=4.655e-13 PD=5.1e-07 PS=1.93e-06
mXSRL/MM57 N_XSRL/SA1_XSRL/MM57_d N_SAEN_XSRL/MM57_g N_DOUT<1>_XSRL/MM57_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13
+ AS=2.4225e-13 PD=1.93e-06 PS=5.1e-07
mXSRL/MM60 N_XSRL/SA1_XSRL/MM60_d N_XSRL/NET0116_XSRL/MM60_g N_VSS_XSRL/MM60_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13
+ AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXSRL/MM61 N_XSRL/NET0116_XSRL/MM61_d N_DOUT_SA<1>_XSRL/MM61_g N_VSS_XSRL/MM61_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13
+ AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXMUX/XI51/MM0 N_BL<9>_XMUX/XI51/MM0_d N_XMUX/NET100_XMUX/XI51/MM0_g
+ N_DL<1>_XMUX/XI51/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI49/MM0 N_BL<10>_XMUX/XI49/MM0_d N_XMUX/NET130_XMUX/XI49/MM0_g
+ N_DL<1>_XMUX/XI49/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSA/MM9 N_XSA/NET012_XSA/MM9_d N_SAEN_XSA/MM9_g N_VSS_XSA/MM9_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXMUX/XI53/MM0 N_BL<11>_XMUX/XI53/MM0_d N_XMUX/NET154_XMUX/XI53/MM0_g
+ N_DL<1>_XMUX/XI53/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI52/MM0 N_BL<12>_XMUX/XI52/MM0_d N_XMUX/NET56_XMUX/XI52/MM0_g
+ N_DL<1>_XMUX/XI52/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI50/MM0 N_BL<13>_XMUX/XI50/MM0_d N_XMUX/NET106_XMUX/XI50/MM0_g
+ N_DL<1>_XMUX/XI50/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI54/MM0 N_BL<14>_XMUX/XI54/MM0_d N_XMUX/NET068_XMUX/XI54/MM0_g
+ N_DL<1>_XMUX/XI54/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSA/MM6 N_XSA/NET016_XSA/MM6_d N_VREF_XSA/MM6_g N_XSA/NET012_XSA/MM6_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.28e-13
+ AS=2.45e-13 PD=5.12e-07 PS=1.48e-06
mXSA/MM3 N_DOUT_SA<1>_XSA/MM3_d N_O1_XSA/MM3_g N_XSA/NET016_XSA/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.28e-13 PD=1.48e-06 PS=5.12e-07
mXMUX/XI48/MM0 N_BL<15>_XMUX/XI48/MM0_d N_XMUX/NET44_XMUX/XI48/MM0_g
+ N_DL<1>_XMUX/XI48/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI2/MM0
+ N_XDFF_TIMING_CONTROL/XI9/XI2/NET41_XDFF_Timing_control/XI9/XI2/MM0_d
+ N_CLK_XDFF_Timing_control/XI9/XI2/MM0_g
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=6e-07 W=1.85e-06 AD=1.0915e-12
+ AS=9.065e-13 PD=3.03e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI2/MM1
+ N_XDFF_TIMING_CONTROL/XI9/XI2/NET37_XDFF_Timing_control/XI9/XI2/MM1_d
+ N_XDFF_TIMING_CONTROL/XI9/XI2/NET41_XDFF_Timing_control/XI9/XI2/MM1_g
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM1_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=6e-07 W=1.85e-06 AD=1.0915e-12
+ AS=9.065e-13 PD=3.03e-06 PS=2.83e-06
mXYDec/XI17/MP N_XYDEC/NET22_XYDec/XI17/MP_d N_Y_SEL_FF<0>_XYDec/XI17/MP_g
+ N_VDD_XYDec/XI17/MP_s N_VDD_XYDec/XI17/MP_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/XI2/MM2
+ N_XDFF_TIMING_CONTROL/XI9/XI2/NET33_XDFF_Timing_control/XI9/XI2/MM2_d
+ N_XDFF_TIMING_CONTROL/XI9/XI2/NET37_XDFF_Timing_control/XI9/XI2/MM2_g
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM2_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=6e-07 W=1.85e-06 AD=1.0915e-12
+ AS=9.065e-13 PD=3.03e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI2/MM3
+ N_XDFF_TIMING_CONTROL/XI9/NET10_XDFF_Timing_control/XI9/XI2/MM3_d
+ N_XDFF_TIMING_CONTROL/XI9/XI2/NET33_XDFF_Timing_control/XI9/XI2/MM3_g
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM3_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=6e-07 W=1.85e-06 AD=1.0915e-12
+ AS=9.065e-13 PD=3.03e-06 PS=2.83e-06
mXYDec/XI18/MP N_XYDEC/NET18_XYDec/XI18/MP_d N_Y_SEL_FF<1>_XYDec/XI18/MP_g
+ N_VDD_XYDec/XI18/MP_s N_VDD_XYDec/XI18/MP_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/MMMb
+ N_XDFF_TIMING_CONTROL/XI9/NET023_XDFF_Timing_control/XI9/MMMb_d
+ N_XDFF_TIMING_CONTROL/XI9/NET10_XDFF_Timing_control/XI9/MMMb_g
+ N_VDD_XDFF_Timing_control/XI9/MMMb_s N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b
+ P_18 L=1e-06 W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXYDec/XI19/MP N_XYDEC/NET14_XYDec/XI19/MP_d N_Y_SEL_FF<2>_XYDec/XI19/MP_g
+ N_VDD_XYDec/XI19/MP_s N_VDD_XYDec/XI19/MP_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI9/MMMd
+ N_XDFF_TIMING_CONTROL/XI9/NET013_XDFF_Timing_control/XI9/MMMd_d
+ N_XDFF_TIMING_CONTROL/XI9/NET023_XDFF_Timing_control/XI9/MMMd_g
+ N_VDD_XDFF_Timing_control/XI9/MMMd_s N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b
+ P_18 L=1e-06 W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI1/XI2/MM0
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI2/NET41_XDFF_Timing_control/XI9/XI1/XI2/MM0_d
+ N_XDFF_TIMING_CONTROL/XI9/NET013_XDFF_Timing_control/XI9/XI1/XI2/MM0_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI2/MM0_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=6e-07 W=1.85e-06 AD=1.0915e-12
+ AS=9.065e-13 PD=3.03e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI2/MM0
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI2/NET41_XDFF_Timing_control/XI9/XI0/XI2/MM0_d
+ N_CLK_XDFF_Timing_control/XI9/XI0/XI2/MM0_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=6e-07 W=1.85e-06
+ AD=1.0915e-12 AS=9.065e-13 PD=3.03e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI1/XI2/MM1
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI2/NET37_XDFF_Timing_control/XI9/XI1/XI2/MM1_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI2/NET41_XDFF_Timing_control/XI9/XI1/XI2/MM1_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI2/MM1_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=6e-07 W=1.85e-06 AD=1.0915e-12
+ AS=9.065e-13 PD=3.03e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI2/MM1
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI2/NET37_XDFF_Timing_control/XI9/XI0/XI2/MM1_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI2/NET41_XDFF_Timing_control/XI9/XI0/XI2/MM1_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM1_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=6e-07 W=1.85e-06
+ AD=1.0915e-12 AS=9.065e-13 PD=3.03e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI1/XI2/MM2
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI2/NET33_XDFF_Timing_control/XI9/XI1/XI2/MM2_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI2/NET37_XDFF_Timing_control/XI9/XI1/XI2/MM2_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI2/MM2_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=6e-07 W=1.85e-06 AD=1.0915e-12
+ AS=9.065e-13 PD=3.03e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI2/MM2
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI2/NET33_XDFF_Timing_control/XI9/XI0/XI2/MM2_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI2/NET37_XDFF_Timing_control/XI9/XI0/XI2/MM2_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM2_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=6e-07 W=1.85e-06
+ AD=1.0915e-12 AS=9.065e-13 PD=3.03e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI1/XI2/MM3
+ N_XDFF_TIMING_CONTROL/XI9/XI1/NET011_XDFF_Timing_control/XI9/XI1/XI2/MM3_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI2/NET33_XDFF_Timing_control/XI9/XI1/XI2/MM3_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI2/MM3_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=6e-07 W=1.85e-06 AD=1.0915e-12
+ AS=9.065e-13 PD=3.03e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI2/MM3
+ N_XDFF_TIMING_CONTROL/XI9/XI0/NET011_XDFF_Timing_control/XI9/XI0/XI2/MM3_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI2/NET33_XDFF_Timing_control/XI9/XI0/XI2/MM3_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM3_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=6e-07 W=1.85e-06
+ AD=1.0915e-12 AS=9.065e-13 PD=3.03e-06 PS=2.83e-06
mXYDec/XI21/MM7 N_Y_SEL<6>_XYDec/XI21/MM7_d N_VDD_XYDec/XI21/MM7_g
+ N_VDD_XYDec/XI21/MM7_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI22/MM7 N_Y_SEL<5>_XYDec/XI22/MM7_d N_VDD_XYDec/XI22/MM7_g
+ N_VDD_XYDec/XI22/MM7_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI25/MM7 N_Y_SEL<2>_XYDec/XI25/MM7_d N_VDD_XYDec/XI25/MM7_g
+ N_VDD_XYDec/XI25/MM7_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI26/MM7 N_Y_SEL<1>_XYDec/XI26/MM7_d N_VDD_XYDec/XI26/MM7_g
+ N_VDD_XYDec/XI26/MM7_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI21/MM4 N_Y_SEL<6>_XYDec/XI21/MM4_d N_Y_SEL_FF<2>_XYDec/XI21/MM4_g
+ N_VDD_XYDec/XI21/MM4_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI22/MM4 N_Y_SEL<5>_XYDec/XI22/MM4_d N_Y_SEL_FF<2>_XYDec/XI22/MM4_g
+ N_VDD_XYDec/XI22/MM4_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI25/MM4 N_Y_SEL<2>_XYDec/XI25/MM4_d N_XYDEC/NET14_XYDec/XI25/MM4_g
+ N_VDD_XYDec/XI25/MM4_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI26/MM4 N_Y_SEL<1>_XYDec/XI26/MM4_d N_XYDEC/NET14_XYDec/XI26/MM4_g
+ N_VDD_XYDec/XI26/MM4_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXDFF_Timing_control/XI9/XI1/XI1/MM0
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET39_XDFF_Timing_control/XI9/XI1/XI1/MM0_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/NET011_XDFF_Timing_control/XI9/XI1/XI1/MM0_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI1/MM0_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=1e-06 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI1/MM0
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET39_XDFF_Timing_control/XI9/XI0/XI1/MM0_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/NET011_XDFF_Timing_control/XI9/XI0/XI1/MM0_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI1/MM0_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=1e-06 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXYDec/XI21/MM5 N_Y_SEL<6>_XYDec/XI21/MM5_d N_Y_SEL_FF<1>_XYDec/XI21/MM5_g
+ N_VDD_XYDec/XI21/MM5_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI22/MM5 N_Y_SEL<5>_XYDec/XI22/MM5_d N_XYDEC/NET18_XYDec/XI22/MM5_g
+ N_VDD_XYDec/XI22/MM5_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI25/MM5 N_Y_SEL<2>_XYDec/XI25/MM5_d N_Y_SEL_FF<1>_XYDec/XI25/MM5_g
+ N_VDD_XYDec/XI25/MM5_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI26/MM5 N_Y_SEL<1>_XYDec/XI26/MM5_d N_XYDEC/NET18_XYDec/XI26/MM5_g
+ N_VDD_XYDec/XI26/MM5_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI21/MM6 N_Y_SEL<6>_XYDec/XI21/MM6_d N_XYDEC/NET22_XYDec/XI21/MM6_g
+ N_VDD_XYDec/XI21/MM6_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI22/MM6 N_Y_SEL<5>_XYDec/XI22/MM6_d N_Y_SEL_FF<0>_XYDec/XI22/MM6_g
+ N_VDD_XYDec/XI22/MM6_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI25/MM6 N_Y_SEL<2>_XYDec/XI25/MM6_d N_XYDEC/NET22_XYDec/XI25/MM6_g
+ N_VDD_XYDec/XI25/MM6_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI26/MM6 N_Y_SEL<1>_XYDec/XI26/MM6_d N_Y_SEL_FF<0>_XYDec/XI26/MM6_g
+ N_VDD_XYDec/XI26/MM6_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI20/MM7 N_Y_SEL<7>_XYDec/XI20/MM7_d N_VDD_XYDec/XI20/MM7_g
+ N_VDD_XYDec/XI20/MM7_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI23/MM7 N_Y_SEL<4>_XYDec/XI23/MM7_d N_VDD_XYDec/XI23/MM7_g
+ N_VDD_XYDec/XI23/MM7_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI24/MM7 N_Y_SEL<3>_XYDec/XI24/MM7_d N_VDD_XYDec/XI24/MM7_g
+ N_VDD_XYDec/XI24/MM7_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI27/MM7 N_Y_SEL<0>_XYDec/XI27/MM7_d N_VDD_XYDec/XI27/MM7_g
+ N_VDD_XYDec/XI27/MM7_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI9/XI1/XI1/MM1
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET15_XDFF_Timing_control/XI9/XI1/XI1/MM1_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET39_XDFF_Timing_control/XI9/XI1/XI1/MM1_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI1/MM1_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=1e-06 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI1/MM1
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET15_XDFF_Timing_control/XI9/XI0/XI1/MM1_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET39_XDFF_Timing_control/XI9/XI0/XI1/MM1_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI1/MM1_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=1e-06 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXYDec/XI20/MM4 N_Y_SEL<7>_XYDec/XI20/MM4_d N_Y_SEL_FF<2>_XYDec/XI20/MM4_g
+ N_VDD_XYDec/XI20/MM4_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI23/MM4 N_Y_SEL<4>_XYDec/XI23/MM4_d N_Y_SEL_FF<2>_XYDec/XI23/MM4_g
+ N_VDD_XYDec/XI23/MM4_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI24/MM4 N_Y_SEL<3>_XYDec/XI24/MM4_d N_XYDEC/NET14_XYDec/XI24/MM4_g
+ N_VDD_XYDec/XI24/MM4_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI27/MM4 N_Y_SEL<0>_XYDec/XI27/MM4_d N_XYDEC/NET14_XYDec/XI27/MM4_g
+ N_VDD_XYDec/XI27/MM4_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI20/MM5 N_Y_SEL<7>_XYDec/XI20/MM5_d N_Y_SEL_FF<1>_XYDec/XI20/MM5_g
+ N_VDD_XYDec/XI20/MM5_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI23/MM5 N_Y_SEL<4>_XYDec/XI23/MM5_d N_XYDEC/NET18_XYDec/XI23/MM5_g
+ N_VDD_XYDec/XI23/MM5_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI24/MM5 N_Y_SEL<3>_XYDec/XI24/MM5_d N_Y_SEL_FF<1>_XYDec/XI24/MM5_g
+ N_VDD_XYDec/XI24/MM5_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI27/MM5 N_Y_SEL<0>_XYDec/XI27/MM5_d N_XYDEC/NET18_XYDec/XI27/MM5_g
+ N_VDD_XYDec/XI27/MM5_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXYDec/XI20/MM6 N_Y_SEL<7>_XYDec/XI20/MM6_d N_Y_SEL_FF<0>_XYDec/XI20/MM6_g
+ N_VDD_XYDec/XI20/MM6_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI23/MM6 N_Y_SEL<4>_XYDec/XI23/MM6_d N_XYDEC/NET22_XYDec/XI23/MM6_g
+ N_VDD_XYDec/XI23/MM6_s N_VDD_XYDec/XI21/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI24/MM6 N_Y_SEL<3>_XYDec/XI24/MM6_d N_Y_SEL_FF<0>_XYDec/XI24/MM6_g
+ N_VDD_XYDec/XI24/MM6_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXYDec/XI27/MM6 N_Y_SEL<0>_XYDec/XI27/MM6_d N_XYDEC/NET22_XYDec/XI27/MM6_g
+ N_VDD_XYDec/XI27/MM6_s N_VDD_XYDec/XI25/MM7_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI9/XI1/XI1/MM2
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET31_XDFF_Timing_control/XI9/XI1/XI1/MM2_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET15_XDFF_Timing_control/XI9/XI1/XI1/MM2_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI1/MM2_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=1e-06 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI1/MM2
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET31_XDFF_Timing_control/XI9/XI0/XI1/MM2_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET15_XDFF_Timing_control/XI9/XI0/XI1/MM2_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI1/MM2_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=1e-06 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/MM0 N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/MM0_d
+ N_CLK_XDFF_Timing_control/MM0_g N_VDD_XDFF_Timing_control/MM0_s
+ N_VDD_XDFF_Timing_control/MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI9/XI1/XI1/MM3
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET27_XDFF_Timing_control/XI9/XI1/XI1/MM3_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET31_XDFF_Timing_control/XI9/XI1/XI1/MM3_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI1/MM3_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=1e-06 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI1/MM3
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET27_XDFF_Timing_control/XI9/XI0/XI1/MM3_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET31_XDFF_Timing_control/XI9/XI0/XI1/MM3_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI1/MM3_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=1e-06 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI1/XI1/MM4
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET046_XDFF_Timing_control/XI9/XI1/XI1/MM4_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET27_XDFF_Timing_control/XI9/XI1/XI1/MM4_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI1/MM4_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=1e-06 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI1/MM4
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET046_XDFF_Timing_control/XI9/XI0/XI1/MM4_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET27_XDFF_Timing_control/XI9/XI0/XI1/MM4_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI1/MM4_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=1e-06 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI1/XI1/MMb
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET038_XDFF_Timing_control/XI9/XI1/XI1/MMb_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET046_XDFF_Timing_control/XI9/XI1/XI1/MMb_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI1/MMb_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=1e-06 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI1/MMb
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET038_XDFF_Timing_control/XI9/XI0/XI1/MMb_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET046_XDFF_Timing_control/XI9/XI0/XI1/MMb_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI1/MMb_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=1e-06 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI1/XI1/MMd
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET034_XDFF_Timing_control/XI9/XI1/XI1/MMd_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET038_XDFF_Timing_control/XI9/XI1/XI1/MMd_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI1/MMd_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=1e-06 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI1/MMd
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET034_XDFF_Timing_control/XI9/XI0/XI1/MMd_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET038_XDFF_Timing_control/XI9/XI0/XI1/MMd_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI1/MMd_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=1e-06 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI1/XI1/MMf
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET030_XDFF_Timing_control/XI9/XI1/XI1/MMf_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET034_XDFF_Timing_control/XI9/XI1/XI1/MMf_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI1/MMf_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=1e-06 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI1/MMf
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET030_XDFF_Timing_control/XI9/XI0/XI1/MMf_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET034_XDFF_Timing_control/XI9/XI0/XI1/MMf_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI1/MMf_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=1e-06 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI1/XI1/MMh
+ N_XDFF_TIMING_CONTROL/XI9/XI1/NET6_XDFF_Timing_control/XI9/XI1/XI1/MMh_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI1/NET030_XDFF_Timing_control/XI9/XI1/XI1/MMh_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI1/MMh_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=1e-06 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI1/MMh
+ N_XDFF_TIMING_CONTROL/XI9/XI0/NET6_XDFF_Timing_control/XI9/XI0/XI1/MMh_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI1/NET030_XDFF_Timing_control/XI9/XI0/XI1/MMh_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI1/MMh_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=1e-06 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI1/XI0/MM0
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI0/NET055_XDFF_Timing_control/XI9/XI1/XI0/MM0_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/NET011_XDFF_Timing_control/XI9/XI1/XI0/MM0_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI0/MM0_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXDFF_Timing_control/XI9/XI0/XI0/MM0
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI0/NET055_XDFF_Timing_control/XI9/XI0/XI0/MM0_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/NET011_XDFF_Timing_control/XI9/XI0/XI0/MM0_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI0/MM0_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXDFF_Timing_control/XI9/XI1/XI0/MM1
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI0/NET055_XDFF_Timing_control/XI9/XI1/XI0/MM1_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/NET6_XDFF_Timing_control/XI9/XI1/XI0/MM1_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI0/MM1_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXDFF_Timing_control/XI9/XI0/XI0/MM1
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI0/NET055_XDFF_Timing_control/XI9/XI0/XI0/MM1_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/NET6_XDFF_Timing_control/XI9/XI0/XI0/MM1_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI0/MM1_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXDFF_Timing_control/XI9/XI1/XI0/MM5
+ N_SAEN_XDFF_Timing_control/XI9/XI1/XI0/MM5_d
+ N_XDFF_TIMING_CONTROL/XI9/XI1/XI0/NET055_XDFF_Timing_control/XI9/XI1/XI0/MM5_g
+ N_VDD_XDFF_Timing_control/XI9/XI1/XI0/MM5_s
+ N_VDD_XDFF_Timing_control/XI9/XI2/MM0_b P_18 L=1.8e-07 W=1.85e-06 AD=9.065e-13
+ AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXDFF_Timing_control/XI9/XI0/XI0/MM5
+ N_WL_EN_XDFF_Timing_control/XI9/XI0/XI0/MM5_d
+ N_XDFF_TIMING_CONTROL/XI9/XI0/XI0/NET055_XDFF_Timing_control/XI9/XI0/XI0/MM5_g
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI0/MM5_s
+ N_VDD_XDFF_Timing_control/XI9/XI0/XI2/MM0_b P_18 L=1.8e-07 W=1.85e-06
+ AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXMUX/XI63/MM0 N_XMUX/NET44_XMUX/XI63/MM0_d N_Y_SEL<7>_XMUX/XI63/MM0_g
+ N_VDD_XMUX/XI63/MM0_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI62/MM0 N_XMUX/NET068_XMUX/XI62/MM0_d N_Y_SEL<6>_XMUX/XI62/MM0_g
+ N_VDD_XMUX/XI62/MM0_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI61/MM0 N_XMUX/NET106_XMUX/XI61/MM0_d N_Y_SEL<5>_XMUX/XI61/MM0_g
+ N_VDD_XMUX/XI61/MM0_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI60/MM0 N_XMUX/NET56_XMUX/XI60/MM0_d N_Y_SEL<4>_XMUX/XI60/MM0_g
+ N_VDD_XMUX/XI60/MM0_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI59/MM0 N_XMUX/NET154_XMUX/XI59/MM0_d N_Y_SEL<3>_XMUX/XI59/MM0_g
+ N_VDD_XMUX/XI59/MM0_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI58/MM0 N_XMUX/NET130_XMUX/XI58/MM0_d N_Y_SEL<2>_XMUX/XI58/MM0_g
+ N_VDD_XMUX/XI58/MM0_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI57/MM0 N_XMUX/NET100_XMUX/XI57/MM0_d N_Y_SEL<1>_XMUX/XI57/MM0_g
+ N_VDD_XMUX/XI57/MM0_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI56/MM0 N_XMUX/NET044_XMUX/XI56/MM0_d N_Y_SEL<0>_XMUX/XI56/MM0_g
+ N_VDD_XMUX/XI56/MM0_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXprech/MM0 N_BL<0>_Xprech/MM0_d N_CLK_Xprech/MM0_g N_VDD_Xprech/MM0_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXprech/MM1 N_BL<1>_Xprech/MM1_d N_CLK_Xprech/MM1_g N_VDD_Xprech/MM1_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXMUX/XI40/MM1 N_DL<0>_XMUX/XI40/MM1_d N_Y_SEL<0>_XMUX/XI40/MM1_g
+ N_BL<0>_XMUX/XI40/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSRL/MM16 N_XSRL/CLKB_XSRL/MM16_d N_SAEN_XSRL/MM16_g N_VDD_XSRL/MM16_s
+ N_VDD_XSRL/MM16_b P_18 L=1.8e-07 W=1.43e-06 AD=7.007e-13 AS=7.007e-13
+ PD=2.41e-06 PS=2.41e-06
mXMUX/XI41/MM1 N_DL<0>_XMUX/XI41/MM1_d N_Y_SEL<1>_XMUX/XI41/MM1_g
+ N_BL<1>_XMUX/XI41/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXprech/MM2 N_BL<2>_Xprech/MM2_d N_CLK_Xprech/MM2_g N_VDD_Xprech/MM2_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXMUX/XI42/MM1 N_DL<0>_XMUX/XI42/MM1_d N_Y_SEL<2>_XMUX/XI42/MM1_g
+ N_BL<2>_XMUX/XI42/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXprech/MM3 N_BL<3>_Xprech/MM3_d N_CLK_Xprech/MM3_g N_VDD_Xprech/MM3_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXSA/MM17 N_O0_XSA/MM17_d N_SAEN_XSA/MM17_g N_VDD_XSA/MM17_s N_VDD_XSA/MM17_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXMUX/XI43/MM1 N_DL<0>_XMUX/XI43/MM1_d N_Y_SEL<3>_XMUX/XI43/MM1_g
+ N_BL<3>_XMUX/XI43/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI44/MM1 N_DL<0>_XMUX/XI44/MM1_d N_Y_SEL<4>_XMUX/XI44/MM1_g
+ N_BL<4>_XMUX/XI44/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSA/MM12 N_O0_XSA/MM12_d N_DOUT_SA<0>_XSA/MM12_g N_VDD_XSA/MM12_s
+ N_VDD_XSA/MM17_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXSRL/MM14 N_QB<0>_XSRL/MM14_d N_DOUT<0>_XSRL/MM14_g N_VDD_XSRL/MM14_s
+ N_VDD_XSRL/MM16_b P_18 L=1.8e-07 W=1.43e-06 AD=7.007e-13 AS=7.007e-13
+ PD=2.41e-06 PS=2.41e-06
mXSRL/MM13 N_XSRL/NET0180_XSRL/MM13_d N_QB<0>_XSRL/MM13_g N_VDD_XSRL/MM13_s
+ N_VDD_XSRL/MM16_b P_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13 AS=4.655e-13
+ PD=1.93e-06 PS=1.93e-06
mXSRL/MM18 N_XSRL/SA0_XSRL/MM18_d N_XSRL/NET088_XSRL/MM18_g N_VDD_XSRL/MM18_s
+ N_VDD_XSRL/MM16_b P_18 L=1.8e-07 W=1.43e-06 AD=7.007e-13 AS=7.007e-13
+ PD=2.41e-06 PS=2.41e-06
mXSRL/MM22 N_XSRL/NET088_XSRL/MM22_d N_DOUT_SA<0>_XSRL/MM22_g N_VDD_XSRL/MM22_s
+ N_VDD_XSRL/MM16_b P_18 L=1.8e-07 W=1.43e-06 AD=7.007e-13 AS=7.007e-13
+ PD=2.41e-06 PS=2.41e-06
mXprech/MM4 N_BL<4>_Xprech/MM4_d N_CLK_Xprech/MM4_g N_VDD_Xprech/MM4_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXSRL/MM40 N_DOUT<0>_XSRL/MM40_d N_SAEN_XSRL/MM40_g N_XSRL/NET0180_XSRL/MM40_s
+ N_VDD_XSRL/MM16_b P_18 L=1.8e-07 W=9.5e-07 AD=2.4225e-13 AS=4.655e-13
+ PD=5.1e-07 PS=1.93e-06
mXSRL/MM17 N_XSRL/SA0_XSRL/MM17_d N_XSRL/CLKB_XSRL/MM17_g N_DOUT<0>_XSRL/MM17_s
+ N_VDD_XSRL/MM16_b P_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13 AS=2.4225e-13
+ PD=1.93e-06 PS=5.1e-07
mXMUX/XI45/MM1 N_DL<0>_XMUX/XI45/MM1_d N_Y_SEL<5>_XMUX/XI45/MM1_g
+ N_BL<5>_XMUX/XI45/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXprech/MM5 N_BL<5>_Xprech/MM5_d N_CLK_Xprech/MM5_g N_VDD_Xprech/MM5_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXMUX/XI46/MM1 N_DL<0>_XMUX/XI46/MM1_d N_Y_SEL<6>_XMUX/XI46/MM1_g
+ N_BL<6>_XMUX/XI46/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSA/MM14 N_DOUT_SA<0>_XSA/MM14_d N_O0_XSA/MM14_g N_VDD_XSA/MM14_s
+ N_VDD_XSA/MM17_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXMUX/XI47/MM1 N_DL<0>_XMUX/XI47/MM1_d N_Y_SEL<7>_XMUX/XI47/MM1_g
+ N_BL<7>_XMUX/XI47/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSA/MM18 N_DOUT_SA<0>_XSA/MM18_d N_SAEN_XSA/MM18_g N_VDD_XSA/MM18_s
+ N_VDD_XSA/MM17_b P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13
+ PD=5.1e-07 PS=1.45e-06
mXprech/MM6 N_BL<6>_Xprech/MM6_d N_CLK_Xprech/MM6_g N_VDD_Xprech/MM6_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXprech/MM7 N_BL<7>_Xprech/MM7_d N_CLK_Xprech/MM7_g N_VDD_Xprech/MM7_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXMUX/XI55/MM1 N_DL<1>_XMUX/XI55/MM1_d N_Y_SEL<0>_XMUX/XI55/MM1_g
+ N_BL<8>_XMUX/XI55/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXprech/MM8 N_BL<8>_Xprech/MM8_d N_CLK_Xprech/MM8_g N_VDD_Xprech/MM8_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXMUX/XI51/MM1 N_DL<1>_XMUX/XI51/MM1_d N_Y_SEL<1>_XMUX/XI51/MM1_g
+ N_BL<9>_XMUX/XI51/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXMUX/XI49/MM1 N_DL<1>_XMUX/XI49/MM1_d N_Y_SEL<2>_XMUX/XI49/MM1_g
+ N_BL<10>_XMUX/XI49/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXprech/MM9 N_BL<9>_Xprech/MM9_d N_CLK_Xprech/MM9_g N_VDD_Xprech/MM9_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXMUX/XI53/MM1 N_DL<1>_XMUX/XI53/MM1_d N_Y_SEL<3>_XMUX/XI53/MM1_g
+ N_BL<11>_XMUX/XI53/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSA/MM7 N_O1_XSA/MM7_d N_SAEN_XSA/MM7_g N_VDD_XSA/MM7_s N_VDD_XSA/MM7_b P_18
+ L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXMUX/XI52/MM1 N_DL<1>_XMUX/XI52/MM1_d N_Y_SEL<4>_XMUX/XI52/MM1_g
+ N_BL<12>_XMUX/XI52/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXprech/MM10 N_BL<10>_Xprech/MM10_d N_CLK_Xprech/MM10_g N_VDD_Xprech/MM10_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXSA/MM2 N_O1_XSA/MM2_d N_DOUT_SA<1>_XSA/MM2_g N_VDD_XSA/MM2_s N_VDD_XSA/MM7_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXMUX/XI50/MM1 N_DL<1>_XMUX/XI50/MM1_d N_Y_SEL<5>_XMUX/XI50/MM1_g
+ N_BL<13>_XMUX/XI50/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXprech/MM11 N_BL<11>_Xprech/MM11_d N_CLK_Xprech/MM11_g N_VDD_Xprech/MM11_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXSRL/MM53 N_QB<1>_XSRL/MM53_d N_DOUT<1>_XSRL/MM53_g N_VDD_XSRL/MM53_s
+ N_VDD_XSRL/MM53_b P_18 L=1.8e-07 W=1.43e-06 AD=7.007e-13 AS=7.007e-13
+ PD=2.41e-06 PS=2.41e-06
mXSRL/MM50 N_DOUT<1>_XSRL/MM50_d N_SAEN_XSRL/MM50_g N_XSRL/NET0178_XSRL/MM50_s
+ N_VDD_XSRL/MM53_b P_18 L=1.8e-07 W=9.5e-07 AD=2.4225e-13 AS=4.655e-13
+ PD=5.1e-07 PS=1.93e-06
mXSRL/MM52 N_XSRL/SA1_XSRL/MM52_d N_XSRL/CLKB_XSRL/MM52_g N_DOUT<1>_XSRL/MM52_s
+ N_VDD_XSRL/MM53_b P_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13 AS=2.4225e-13
+ PD=1.93e-06 PS=5.1e-07
mXSRL/MM58 N_XSRL/SA1_XSRL/MM58_d N_XSRL/NET0116_XSRL/MM58_g N_VDD_XSRL/MM58_s
+ N_VDD_XSRL/MM53_b P_18 L=1.8e-07 W=1.43e-06 AD=7.007e-13 AS=7.007e-13
+ PD=2.41e-06 PS=2.41e-06
mXSRL/MM59 N_XSRL/NET0116_XSRL/MM59_d N_DOUT_SA<1>_XSRL/MM59_g N_VDD_XSRL/MM59_s
+ N_VDD_XSRL/MM53_b P_18 L=1.8e-07 W=1.43e-06 AD=7.007e-13 AS=7.007e-13
+ PD=2.41e-06 PS=2.41e-06
mXMUX/XI54/MM1 N_DL<1>_XMUX/XI54/MM1_d N_Y_SEL<6>_XMUX/XI54/MM1_g
+ N_BL<14>_XMUX/XI54/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSRL/MM51 N_XSRL/NET0178_XSRL/MM51_d N_QB<1>_XSRL/MM51_g N_VDD_XSRL/MM51_s
+ N_VDD_XSRL/MM53_b P_18 L=1.8e-07 W=9.5e-07 AD=4.655e-13 AS=4.655e-13
+ PD=1.93e-06 PS=1.93e-06
mXMUX/XI48/MM1 N_DL<1>_XMUX/XI48/MM1_d N_Y_SEL<7>_XMUX/XI48/MM1_g
+ N_BL<15>_XMUX/XI48/MM1_s N_VDD_XMUX/XI63/MM0_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXSA/MM4 N_DOUT_SA<1>_XSA/MM4_d N_O1_XSA/MM4_g N_VDD_XSA/MM4_s N_VDD_XSA/MM7_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXprech/MM12 N_BL<12>_Xprech/MM12_d N_CLK_Xprech/MM12_g N_VDD_Xprech/MM12_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXSA/MM8 N_DOUT_SA<1>_XSA/MM8_d N_SAEN_XSA/MM8_g N_VDD_XSA/MM8_s N_VDD_XSA/MM7_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXprech/MM13 N_BL<13>_Xprech/MM13_d N_CLK_Xprech/MM13_g N_VDD_Xprech/MM13_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXprech/MM14 N_BL<14>_Xprech/MM14_d N_CLK_Xprech/MM14_g N_VDD_Xprech/MM14_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXprech/MM15 N_BL<15>_Xprech/MM15_d N_CLK_Xprech/MM15_g N_VDD_Xprech/MM15_s
+ N_VDD_Xprech/MM0_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=1.1985e-13
+ PD=1.45e-06 PS=5.1e-07
mXDFF_Timing_control/XI3/MM0
+ N_XDFF_TIMING_CONTROL/XI3/NET92_XDFF_Timing_control/XI3/MM0_d
+ N_A<2>_XDFF_Timing_control/XI3/MM0_g N_VSS_XDFF_Timing_control/XI3/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI3/MM10
+ N_XDFF_TIMING_CONTROL/XI3/NET92_XDFF_Timing_control/XI3/MM10_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI3/MM10_g
+ N_XDFF_TIMING_CONTROL/XI3/NET75_XDFF_Timing_control/XI3/MM10_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI3/MM3
+ N_XDFF_TIMING_CONTROL/XI3/NET22_XDFF_Timing_control/XI3/MM3_d
+ N_XDFF_TIMING_CONTROL/XI3/NET75_XDFF_Timing_control/XI3/MM3_g
+ N_VSS_XDFF_Timing_control/XI3/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI3/MM16
+ N_XDFF_TIMING_CONTROL/XI3/NET75_XDFF_Timing_control/XI3/MM16_d
+ N_XDFF_TIMING_CONTROL/XI3/NET22_XDFF_Timing_control/XI3/MM16_g
+ N_XDFF_TIMING_CONTROL/XI3/NET60_XDFF_Timing_control/XI3/MM16_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI3/MM20
+ N_XDFF_TIMING_CONTROL/XI3/NET60_XDFF_Timing_control/XI3/MM20_d
+ N_CLK_XDFF_Timing_control/XI3/MM20_g N_VSS_XDFF_Timing_control/XI3/MM20_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI3/MM13
+ N_XDFF_TIMING_CONTROL/XI3/NET22_XDFF_Timing_control/XI3/MM13_d
+ N_CLK_XDFF_Timing_control/XI3/MM13_g
+ N_XDFF_TIMING_CONTROL/XI3/NET71_XDFF_Timing_control/XI3/MM13_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI3/MM4
+ N_XDFF_TIMING_CONTROL/XI3/NET10_XDFF_Timing_control/XI3/MM4_d
+ N_XDFF_TIMING_CONTROL/XI3/NET71_XDFF_Timing_control/XI3/MM4_g
+ N_VSS_XDFF_Timing_control/XI3/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI3/MM24
+ N_XDFF_TIMING_CONTROL/XI3/NET71_XDFF_Timing_control/XI3/MM24_d
+ N_XDFF_TIMING_CONTROL/XI3/NET10_XDFF_Timing_control/XI3/MM24_g
+ N_XDFF_TIMING_CONTROL/XI3/NET56_XDFF_Timing_control/XI3/MM24_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI3/MM21
+ N_XDFF_TIMING_CONTROL/XI3/NET56_XDFF_Timing_control/XI3/MM21_d
+ N_CLK_XDFF_Timing_control/XI3/MM21_g N_VSS_XDFF_Timing_control/XI3/MM21_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI3/MM9 N_X_SEL_FF<2>_XDFF_Timing_control/XI3/MM9_d
+ N_XDFF_TIMING_CONTROL/XI3/NET10_XDFF_Timing_control/XI3/MM9_g
+ N_VSS_XDFF_Timing_control/XI3/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI3/MM7 N_NOTUSED2_XDFF_Timing_control/XI3/MM7_d
+ N_XDFF_TIMING_CONTROL/XI3/NET71_XDFF_Timing_control/XI3/MM7_g
+ N_VSS_XDFF_Timing_control/XI3/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI3/MM1
+ N_XDFF_TIMING_CONTROL/XI3/NET92_XDFF_Timing_control/XI3/MM1_d
+ N_A<2>_XDFF_Timing_control/XI3/MM1_g N_VDD_XDFF_Timing_control/XI3/MM1_s
+ N_VDD_XDFF_Timing_control/XI3/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI3/MM12
+ N_XDFF_TIMING_CONTROL/XI3/NET92_XDFF_Timing_control/XI3/MM12_d
+ N_CLK_XDFF_Timing_control/XI3/MM12_g
+ N_XDFF_TIMING_CONTROL/XI3/NET75_XDFF_Timing_control/XI3/MM12_s
+ N_VDD_XDFF_Timing_control/XI3/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI3/MM2
+ N_XDFF_TIMING_CONTROL/XI3/NET22_XDFF_Timing_control/XI3/MM2_d
+ N_XDFF_TIMING_CONTROL/XI3/NET75_XDFF_Timing_control/XI3/MM2_g
+ N_VDD_XDFF_Timing_control/XI3/MM2_s N_VDD_XDFF_Timing_control/XI3/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI3/MM15
+ N_XDFF_TIMING_CONTROL/XI3/NET75_XDFF_Timing_control/XI3/MM15_d
+ N_XDFF_TIMING_CONTROL/XI3/NET22_XDFF_Timing_control/XI3/MM15_g
+ N_XDFF_TIMING_CONTROL/XI3/NET23_XDFF_Timing_control/XI3/MM15_s
+ N_VDD_XDFF_Timing_control/XI3/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI3/MM19
+ N_XDFF_TIMING_CONTROL/XI3/NET23_XDFF_Timing_control/XI3/MM19_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI3/MM19_g
+ N_VDD_XDFF_Timing_control/XI3/MM19_s N_VDD_XDFF_Timing_control/XI3/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI3/MM11
+ N_XDFF_TIMING_CONTROL/XI3/NET22_XDFF_Timing_control/XI3/MM11_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI3/MM11_g
+ N_XDFF_TIMING_CONTROL/XI3/NET71_XDFF_Timing_control/XI3/MM11_s
+ N_VDD_XDFF_Timing_control/XI3/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI3/MM5
+ N_XDFF_TIMING_CONTROL/XI3/NET10_XDFF_Timing_control/XI3/MM5_d
+ N_XDFF_TIMING_CONTROL/XI3/NET71_XDFF_Timing_control/XI3/MM5_g
+ N_VDD_XDFF_Timing_control/XI3/MM5_s N_VDD_XDFF_Timing_control/XI3/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI3/MM23
+ N_XDFF_TIMING_CONTROL/XI3/NET71_XDFF_Timing_control/XI3/MM23_d
+ N_XDFF_TIMING_CONTROL/XI3/NET10_XDFF_Timing_control/XI3/MM23_g
+ N_XDFF_TIMING_CONTROL/XI3/NET12_XDFF_Timing_control/XI3/MM23_s
+ N_VDD_XDFF_Timing_control/XI3/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI3/MM22
+ N_XDFF_TIMING_CONTROL/XI3/NET12_XDFF_Timing_control/XI3/MM22_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI3/MM22_g
+ N_VDD_XDFF_Timing_control/XI3/MM22_s N_VDD_XDFF_Timing_control/XI3/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI3/MM8 N_X_SEL_FF<2>_XDFF_Timing_control/XI3/MM8_d
+ N_XDFF_TIMING_CONTROL/XI3/NET10_XDFF_Timing_control/XI3/MM8_g
+ N_VDD_XDFF_Timing_control/XI3/MM8_s N_VDD_XDFF_Timing_control/XI3/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI3/MM6 N_NOTUSED2_XDFF_Timing_control/XI3/MM6_d
+ N_XDFF_TIMING_CONTROL/XI3/NET71_XDFF_Timing_control/XI3/MM6_g
+ N_VDD_XDFF_Timing_control/XI3/MM6_s N_VDD_XDFF_Timing_control/XI3/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI6/MM0
+ N_XDFF_TIMING_CONTROL/XI6/NET92_XDFF_Timing_control/XI6/MM0_d
+ N_A<5>_XDFF_Timing_control/XI6/MM0_g N_VSS_XDFF_Timing_control/XI6/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI6/MM10
+ N_XDFF_TIMING_CONTROL/XI6/NET92_XDFF_Timing_control/XI6/MM10_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI6/MM10_g
+ N_XDFF_TIMING_CONTROL/XI6/NET75_XDFF_Timing_control/XI6/MM10_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI6/MM3
+ N_XDFF_TIMING_CONTROL/XI6/NET22_XDFF_Timing_control/XI6/MM3_d
+ N_XDFF_TIMING_CONTROL/XI6/NET75_XDFF_Timing_control/XI6/MM3_g
+ N_VSS_XDFF_Timing_control/XI6/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI6/MM16
+ N_XDFF_TIMING_CONTROL/XI6/NET75_XDFF_Timing_control/XI6/MM16_d
+ N_XDFF_TIMING_CONTROL/XI6/NET22_XDFF_Timing_control/XI6/MM16_g
+ N_XDFF_TIMING_CONTROL/XI6/NET60_XDFF_Timing_control/XI6/MM16_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI6/MM20
+ N_XDFF_TIMING_CONTROL/XI6/NET60_XDFF_Timing_control/XI6/MM20_d
+ N_CLK_XDFF_Timing_control/XI6/MM20_g N_VSS_XDFF_Timing_control/XI6/MM20_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI6/MM13
+ N_XDFF_TIMING_CONTROL/XI6/NET22_XDFF_Timing_control/XI6/MM13_d
+ N_CLK_XDFF_Timing_control/XI6/MM13_g
+ N_XDFF_TIMING_CONTROL/XI6/NET71_XDFF_Timing_control/XI6/MM13_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI6/MM4
+ N_XDFF_TIMING_CONTROL/XI6/NET10_XDFF_Timing_control/XI6/MM4_d
+ N_XDFF_TIMING_CONTROL/XI6/NET71_XDFF_Timing_control/XI6/MM4_g
+ N_VSS_XDFF_Timing_control/XI6/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI6/MM24
+ N_XDFF_TIMING_CONTROL/XI6/NET71_XDFF_Timing_control/XI6/MM24_d
+ N_XDFF_TIMING_CONTROL/XI6/NET10_XDFF_Timing_control/XI6/MM24_g
+ N_XDFF_TIMING_CONTROL/XI6/NET56_XDFF_Timing_control/XI6/MM24_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI6/MM21
+ N_XDFF_TIMING_CONTROL/XI6/NET56_XDFF_Timing_control/XI6/MM21_d
+ N_CLK_XDFF_Timing_control/XI6/MM21_g N_VSS_XDFF_Timing_control/XI6/MM21_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI6/MM9 N_X_SEL_FF<5>_XDFF_Timing_control/XI6/MM9_d
+ N_XDFF_TIMING_CONTROL/XI6/NET10_XDFF_Timing_control/XI6/MM9_g
+ N_VSS_XDFF_Timing_control/XI6/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI6/MM7 N_NOTUSED5_XDFF_Timing_control/XI6/MM7_d
+ N_XDFF_TIMING_CONTROL/XI6/NET71_XDFF_Timing_control/XI6/MM7_g
+ N_VSS_XDFF_Timing_control/XI6/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI6/MM1
+ N_XDFF_TIMING_CONTROL/XI6/NET92_XDFF_Timing_control/XI6/MM1_d
+ N_A<5>_XDFF_Timing_control/XI6/MM1_g N_VDD_XDFF_Timing_control/XI6/MM1_s
+ N_VDD_XDFF_Timing_control/XI6/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI6/MM12
+ N_XDFF_TIMING_CONTROL/XI6/NET92_XDFF_Timing_control/XI6/MM12_d
+ N_CLK_XDFF_Timing_control/XI6/MM12_g
+ N_XDFF_TIMING_CONTROL/XI6/NET75_XDFF_Timing_control/XI6/MM12_s
+ N_VDD_XDFF_Timing_control/XI6/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI6/MM2
+ N_XDFF_TIMING_CONTROL/XI6/NET22_XDFF_Timing_control/XI6/MM2_d
+ N_XDFF_TIMING_CONTROL/XI6/NET75_XDFF_Timing_control/XI6/MM2_g
+ N_VDD_XDFF_Timing_control/XI6/MM2_s N_VDD_XDFF_Timing_control/XI6/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI6/MM15
+ N_XDFF_TIMING_CONTROL/XI6/NET75_XDFF_Timing_control/XI6/MM15_d
+ N_XDFF_TIMING_CONTROL/XI6/NET22_XDFF_Timing_control/XI6/MM15_g
+ N_XDFF_TIMING_CONTROL/XI6/NET23_XDFF_Timing_control/XI6/MM15_s
+ N_VDD_XDFF_Timing_control/XI6/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI6/MM19
+ N_XDFF_TIMING_CONTROL/XI6/NET23_XDFF_Timing_control/XI6/MM19_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI6/MM19_g
+ N_VDD_XDFF_Timing_control/XI6/MM19_s N_VDD_XDFF_Timing_control/XI6/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI6/MM11
+ N_XDFF_TIMING_CONTROL/XI6/NET22_XDFF_Timing_control/XI6/MM11_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI6/MM11_g
+ N_XDFF_TIMING_CONTROL/XI6/NET71_XDFF_Timing_control/XI6/MM11_s
+ N_VDD_XDFF_Timing_control/XI6/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI6/MM5
+ N_XDFF_TIMING_CONTROL/XI6/NET10_XDFF_Timing_control/XI6/MM5_d
+ N_XDFF_TIMING_CONTROL/XI6/NET71_XDFF_Timing_control/XI6/MM5_g
+ N_VDD_XDFF_Timing_control/XI6/MM5_s N_VDD_XDFF_Timing_control/XI6/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI6/MM23
+ N_XDFF_TIMING_CONTROL/XI6/NET71_XDFF_Timing_control/XI6/MM23_d
+ N_XDFF_TIMING_CONTROL/XI6/NET10_XDFF_Timing_control/XI6/MM23_g
+ N_XDFF_TIMING_CONTROL/XI6/NET12_XDFF_Timing_control/XI6/MM23_s
+ N_VDD_XDFF_Timing_control/XI6/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI6/MM22
+ N_XDFF_TIMING_CONTROL/XI6/NET12_XDFF_Timing_control/XI6/MM22_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI6/MM22_g
+ N_VDD_XDFF_Timing_control/XI6/MM22_s N_VDD_XDFF_Timing_control/XI6/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI6/MM8 N_X_SEL_FF<5>_XDFF_Timing_control/XI6/MM8_d
+ N_XDFF_TIMING_CONTROL/XI6/NET10_XDFF_Timing_control/XI6/MM8_g
+ N_VDD_XDFF_Timing_control/XI6/MM8_s N_VDD_XDFF_Timing_control/XI6/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI6/MM6 N_NOTUSED5_XDFF_Timing_control/XI6/MM6_d
+ N_XDFF_TIMING_CONTROL/XI6/NET71_XDFF_Timing_control/XI6/MM6_g
+ N_VDD_XDFF_Timing_control/XI6/MM6_s N_VDD_XDFF_Timing_control/XI6/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI1/MM0
+ N_XDFF_TIMING_CONTROL/XI1/NET92_XDFF_Timing_control/XI1/MM0_d
+ N_A<6>_XDFF_Timing_control/XI1/MM0_g N_VSS_XDFF_Timing_control/XI1/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI1/MM10
+ N_XDFF_TIMING_CONTROL/XI1/NET92_XDFF_Timing_control/XI1/MM10_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI1/MM10_g
+ N_XDFF_TIMING_CONTROL/XI1/NET75_XDFF_Timing_control/XI1/MM10_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI1/MM3
+ N_XDFF_TIMING_CONTROL/XI1/NET22_XDFF_Timing_control/XI1/MM3_d
+ N_XDFF_TIMING_CONTROL/XI1/NET75_XDFF_Timing_control/XI1/MM3_g
+ N_VSS_XDFF_Timing_control/XI1/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI1/MM16
+ N_XDFF_TIMING_CONTROL/XI1/NET75_XDFF_Timing_control/XI1/MM16_d
+ N_XDFF_TIMING_CONTROL/XI1/NET22_XDFF_Timing_control/XI1/MM16_g
+ N_XDFF_TIMING_CONTROL/XI1/NET60_XDFF_Timing_control/XI1/MM16_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI1/MM20
+ N_XDFF_TIMING_CONTROL/XI1/NET60_XDFF_Timing_control/XI1/MM20_d
+ N_CLK_XDFF_Timing_control/XI1/MM20_g N_VSS_XDFF_Timing_control/XI1/MM20_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI1/MM13
+ N_XDFF_TIMING_CONTROL/XI1/NET22_XDFF_Timing_control/XI1/MM13_d
+ N_CLK_XDFF_Timing_control/XI1/MM13_g
+ N_XDFF_TIMING_CONTROL/XI1/NET71_XDFF_Timing_control/XI1/MM13_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI1/MM4
+ N_XDFF_TIMING_CONTROL/XI1/NET10_XDFF_Timing_control/XI1/MM4_d
+ N_XDFF_TIMING_CONTROL/XI1/NET71_XDFF_Timing_control/XI1/MM4_g
+ N_VSS_XDFF_Timing_control/XI1/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI1/MM24
+ N_XDFF_TIMING_CONTROL/XI1/NET71_XDFF_Timing_control/XI1/MM24_d
+ N_XDFF_TIMING_CONTROL/XI1/NET10_XDFF_Timing_control/XI1/MM24_g
+ N_XDFF_TIMING_CONTROL/XI1/NET56_XDFF_Timing_control/XI1/MM24_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI1/MM21
+ N_XDFF_TIMING_CONTROL/XI1/NET56_XDFF_Timing_control/XI1/MM21_d
+ N_CLK_XDFF_Timing_control/XI1/MM21_g N_VSS_XDFF_Timing_control/XI1/MM21_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI1/MM9 N_Y_SEL_FF<0>_XDFF_Timing_control/XI1/MM9_d
+ N_XDFF_TIMING_CONTROL/XI1/NET10_XDFF_Timing_control/XI1/MM9_g
+ N_VSS_XDFF_Timing_control/XI1/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI1/MM7 N_NOTUSED6_XDFF_Timing_control/XI1/MM7_d
+ N_XDFF_TIMING_CONTROL/XI1/NET71_XDFF_Timing_control/XI1/MM7_g
+ N_VSS_XDFF_Timing_control/XI1/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI1/MM1
+ N_XDFF_TIMING_CONTROL/XI1/NET92_XDFF_Timing_control/XI1/MM1_d
+ N_A<6>_XDFF_Timing_control/XI1/MM1_g N_VDD_XDFF_Timing_control/XI1/MM1_s
+ N_VDD_XDFF_Timing_control/XI1/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI1/MM12
+ N_XDFF_TIMING_CONTROL/XI1/NET92_XDFF_Timing_control/XI1/MM12_d
+ N_CLK_XDFF_Timing_control/XI1/MM12_g
+ N_XDFF_TIMING_CONTROL/XI1/NET75_XDFF_Timing_control/XI1/MM12_s
+ N_VDD_XDFF_Timing_control/XI1/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI1/MM2
+ N_XDFF_TIMING_CONTROL/XI1/NET22_XDFF_Timing_control/XI1/MM2_d
+ N_XDFF_TIMING_CONTROL/XI1/NET75_XDFF_Timing_control/XI1/MM2_g
+ N_VDD_XDFF_Timing_control/XI1/MM2_s N_VDD_XDFF_Timing_control/XI1/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI1/MM15
+ N_XDFF_TIMING_CONTROL/XI1/NET75_XDFF_Timing_control/XI1/MM15_d
+ N_XDFF_TIMING_CONTROL/XI1/NET22_XDFF_Timing_control/XI1/MM15_g
+ N_XDFF_TIMING_CONTROL/XI1/NET23_XDFF_Timing_control/XI1/MM15_s
+ N_VDD_XDFF_Timing_control/XI1/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI1/MM19
+ N_XDFF_TIMING_CONTROL/XI1/NET23_XDFF_Timing_control/XI1/MM19_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI1/MM19_g
+ N_VDD_XDFF_Timing_control/XI1/MM19_s N_VDD_XDFF_Timing_control/XI1/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI1/MM11
+ N_XDFF_TIMING_CONTROL/XI1/NET22_XDFF_Timing_control/XI1/MM11_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI1/MM11_g
+ N_XDFF_TIMING_CONTROL/XI1/NET71_XDFF_Timing_control/XI1/MM11_s
+ N_VDD_XDFF_Timing_control/XI1/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI1/MM5
+ N_XDFF_TIMING_CONTROL/XI1/NET10_XDFF_Timing_control/XI1/MM5_d
+ N_XDFF_TIMING_CONTROL/XI1/NET71_XDFF_Timing_control/XI1/MM5_g
+ N_VDD_XDFF_Timing_control/XI1/MM5_s N_VDD_XDFF_Timing_control/XI1/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI1/MM23
+ N_XDFF_TIMING_CONTROL/XI1/NET71_XDFF_Timing_control/XI1/MM23_d
+ N_XDFF_TIMING_CONTROL/XI1/NET10_XDFF_Timing_control/XI1/MM23_g
+ N_XDFF_TIMING_CONTROL/XI1/NET12_XDFF_Timing_control/XI1/MM23_s
+ N_VDD_XDFF_Timing_control/XI1/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI1/MM22
+ N_XDFF_TIMING_CONTROL/XI1/NET12_XDFF_Timing_control/XI1/MM22_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI1/MM22_g
+ N_VDD_XDFF_Timing_control/XI1/MM22_s N_VDD_XDFF_Timing_control/XI1/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI1/MM8 N_Y_SEL_FF<0>_XDFF_Timing_control/XI1/MM8_d
+ N_XDFF_TIMING_CONTROL/XI1/NET10_XDFF_Timing_control/XI1/MM8_g
+ N_VDD_XDFF_Timing_control/XI1/MM8_s N_VDD_XDFF_Timing_control/XI1/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI1/MM6 N_NOTUSED6_XDFF_Timing_control/XI1/MM6_d
+ N_XDFF_TIMING_CONTROL/XI1/NET71_XDFF_Timing_control/XI1/MM6_g
+ N_VDD_XDFF_Timing_control/XI1/MM6_s N_VDD_XDFF_Timing_control/XI1/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI0/MM0
+ N_XDFF_TIMING_CONTROL/XI0/NET92_XDFF_Timing_control/XI0/MM0_d
+ N_A<7>_XDFF_Timing_control/XI0/MM0_g N_VSS_XDFF_Timing_control/XI0/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI0/MM10
+ N_XDFF_TIMING_CONTROL/XI0/NET92_XDFF_Timing_control/XI0/MM10_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI0/MM10_g
+ N_XDFF_TIMING_CONTROL/XI0/NET75_XDFF_Timing_control/XI0/MM10_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI0/MM3
+ N_XDFF_TIMING_CONTROL/XI0/NET22_XDFF_Timing_control/XI0/MM3_d
+ N_XDFF_TIMING_CONTROL/XI0/NET75_XDFF_Timing_control/XI0/MM3_g
+ N_VSS_XDFF_Timing_control/XI0/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI0/MM16
+ N_XDFF_TIMING_CONTROL/XI0/NET75_XDFF_Timing_control/XI0/MM16_d
+ N_XDFF_TIMING_CONTROL/XI0/NET22_XDFF_Timing_control/XI0/MM16_g
+ N_XDFF_TIMING_CONTROL/XI0/NET60_XDFF_Timing_control/XI0/MM16_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI0/MM20
+ N_XDFF_TIMING_CONTROL/XI0/NET60_XDFF_Timing_control/XI0/MM20_d
+ N_CLK_XDFF_Timing_control/XI0/MM20_g N_VSS_XDFF_Timing_control/XI0/MM20_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI0/MM13
+ N_XDFF_TIMING_CONTROL/XI0/NET22_XDFF_Timing_control/XI0/MM13_d
+ N_CLK_XDFF_Timing_control/XI0/MM13_g
+ N_XDFF_TIMING_CONTROL/XI0/NET71_XDFF_Timing_control/XI0/MM13_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI0/MM4
+ N_XDFF_TIMING_CONTROL/XI0/NET10_XDFF_Timing_control/XI0/MM4_d
+ N_XDFF_TIMING_CONTROL/XI0/NET71_XDFF_Timing_control/XI0/MM4_g
+ N_VSS_XDFF_Timing_control/XI0/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI0/MM24
+ N_XDFF_TIMING_CONTROL/XI0/NET71_XDFF_Timing_control/XI0/MM24_d
+ N_XDFF_TIMING_CONTROL/XI0/NET10_XDFF_Timing_control/XI0/MM24_g
+ N_XDFF_TIMING_CONTROL/XI0/NET56_XDFF_Timing_control/XI0/MM24_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI0/MM21
+ N_XDFF_TIMING_CONTROL/XI0/NET56_XDFF_Timing_control/XI0/MM21_d
+ N_CLK_XDFF_Timing_control/XI0/MM21_g N_VSS_XDFF_Timing_control/XI0/MM21_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI0/MM9 N_Y_SEL_FF<1>_XDFF_Timing_control/XI0/MM9_d
+ N_XDFF_TIMING_CONTROL/XI0/NET10_XDFF_Timing_control/XI0/MM9_g
+ N_VSS_XDFF_Timing_control/XI0/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI0/MM7 N_NOTUSED7_XDFF_Timing_control/XI0/MM7_d
+ N_XDFF_TIMING_CONTROL/XI0/NET71_XDFF_Timing_control/XI0/MM7_g
+ N_VSS_XDFF_Timing_control/XI0/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI0/MM1
+ N_XDFF_TIMING_CONTROL/XI0/NET92_XDFF_Timing_control/XI0/MM1_d
+ N_A<7>_XDFF_Timing_control/XI0/MM1_g N_VDD_XDFF_Timing_control/XI0/MM1_s
+ N_VDD_XDFF_Timing_control/XI0/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI0/MM12
+ N_XDFF_TIMING_CONTROL/XI0/NET92_XDFF_Timing_control/XI0/MM12_d
+ N_CLK_XDFF_Timing_control/XI0/MM12_g
+ N_XDFF_TIMING_CONTROL/XI0/NET75_XDFF_Timing_control/XI0/MM12_s
+ N_VDD_XDFF_Timing_control/XI0/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI0/MM2
+ N_XDFF_TIMING_CONTROL/XI0/NET22_XDFF_Timing_control/XI0/MM2_d
+ N_XDFF_TIMING_CONTROL/XI0/NET75_XDFF_Timing_control/XI0/MM2_g
+ N_VDD_XDFF_Timing_control/XI0/MM2_s N_VDD_XDFF_Timing_control/XI0/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI0/MM15
+ N_XDFF_TIMING_CONTROL/XI0/NET75_XDFF_Timing_control/XI0/MM15_d
+ N_XDFF_TIMING_CONTROL/XI0/NET22_XDFF_Timing_control/XI0/MM15_g
+ N_XDFF_TIMING_CONTROL/XI0/NET23_XDFF_Timing_control/XI0/MM15_s
+ N_VDD_XDFF_Timing_control/XI0/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI0/MM19
+ N_XDFF_TIMING_CONTROL/XI0/NET23_XDFF_Timing_control/XI0/MM19_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI0/MM19_g
+ N_VDD_XDFF_Timing_control/XI0/MM19_s N_VDD_XDFF_Timing_control/XI0/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI0/MM11
+ N_XDFF_TIMING_CONTROL/XI0/NET22_XDFF_Timing_control/XI0/MM11_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI0/MM11_g
+ N_XDFF_TIMING_CONTROL/XI0/NET71_XDFF_Timing_control/XI0/MM11_s
+ N_VDD_XDFF_Timing_control/XI0/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI0/MM5
+ N_XDFF_TIMING_CONTROL/XI0/NET10_XDFF_Timing_control/XI0/MM5_d
+ N_XDFF_TIMING_CONTROL/XI0/NET71_XDFF_Timing_control/XI0/MM5_g
+ N_VDD_XDFF_Timing_control/XI0/MM5_s N_VDD_XDFF_Timing_control/XI0/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI0/MM23
+ N_XDFF_TIMING_CONTROL/XI0/NET71_XDFF_Timing_control/XI0/MM23_d
+ N_XDFF_TIMING_CONTROL/XI0/NET10_XDFF_Timing_control/XI0/MM23_g
+ N_XDFF_TIMING_CONTROL/XI0/NET12_XDFF_Timing_control/XI0/MM23_s
+ N_VDD_XDFF_Timing_control/XI0/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI0/MM22
+ N_XDFF_TIMING_CONTROL/XI0/NET12_XDFF_Timing_control/XI0/MM22_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI0/MM22_g
+ N_VDD_XDFF_Timing_control/XI0/MM22_s N_VDD_XDFF_Timing_control/XI0/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI0/MM8 N_Y_SEL_FF<1>_XDFF_Timing_control/XI0/MM8_d
+ N_XDFF_TIMING_CONTROL/XI0/NET10_XDFF_Timing_control/XI0/MM8_g
+ N_VDD_XDFF_Timing_control/XI0/MM8_s N_VDD_XDFF_Timing_control/XI0/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI0/MM6 N_NOTUSED7_XDFF_Timing_control/XI0/MM6_d
+ N_XDFF_TIMING_CONTROL/XI0/NET71_XDFF_Timing_control/XI0/MM6_g
+ N_VDD_XDFF_Timing_control/XI0/MM6_s N_VDD_XDFF_Timing_control/XI0/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI8/MM0
+ N_XDFF_TIMING_CONTROL/XI8/NET92_XDFF_Timing_control/XI8/MM0_d
+ N_A<8>_XDFF_Timing_control/XI8/MM0_g N_VSS_XDFF_Timing_control/XI8/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI8/MM10
+ N_XDFF_TIMING_CONTROL/XI8/NET92_XDFF_Timing_control/XI8/MM10_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI8/MM10_g
+ N_XDFF_TIMING_CONTROL/XI8/NET75_XDFF_Timing_control/XI8/MM10_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI8/MM3
+ N_XDFF_TIMING_CONTROL/XI8/NET22_XDFF_Timing_control/XI8/MM3_d
+ N_XDFF_TIMING_CONTROL/XI8/NET75_XDFF_Timing_control/XI8/MM3_g
+ N_VSS_XDFF_Timing_control/XI8/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI8/MM16
+ N_XDFF_TIMING_CONTROL/XI8/NET75_XDFF_Timing_control/XI8/MM16_d
+ N_XDFF_TIMING_CONTROL/XI8/NET22_XDFF_Timing_control/XI8/MM16_g
+ N_XDFF_TIMING_CONTROL/XI8/NET60_XDFF_Timing_control/XI8/MM16_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI8/MM20
+ N_XDFF_TIMING_CONTROL/XI8/NET60_XDFF_Timing_control/XI8/MM20_d
+ N_CLK_XDFF_Timing_control/XI8/MM20_g N_VSS_XDFF_Timing_control/XI8/MM20_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI8/MM13
+ N_XDFF_TIMING_CONTROL/XI8/NET22_XDFF_Timing_control/XI8/MM13_d
+ N_CLK_XDFF_Timing_control/XI8/MM13_g
+ N_XDFF_TIMING_CONTROL/XI8/NET71_XDFF_Timing_control/XI8/MM13_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI8/MM4
+ N_XDFF_TIMING_CONTROL/XI8/NET10_XDFF_Timing_control/XI8/MM4_d
+ N_XDFF_TIMING_CONTROL/XI8/NET71_XDFF_Timing_control/XI8/MM4_g
+ N_VSS_XDFF_Timing_control/XI8/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI8/MM24
+ N_XDFF_TIMING_CONTROL/XI8/NET71_XDFF_Timing_control/XI8/MM24_d
+ N_XDFF_TIMING_CONTROL/XI8/NET10_XDFF_Timing_control/XI8/MM24_g
+ N_XDFF_TIMING_CONTROL/XI8/NET56_XDFF_Timing_control/XI8/MM24_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI8/MM21
+ N_XDFF_TIMING_CONTROL/XI8/NET56_XDFF_Timing_control/XI8/MM21_d
+ N_CLK_XDFF_Timing_control/XI8/MM21_g N_VSS_XDFF_Timing_control/XI8/MM21_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI8/MM9 N_Y_SEL_FF<2>_XDFF_Timing_control/XI8/MM9_d
+ N_XDFF_TIMING_CONTROL/XI8/NET10_XDFF_Timing_control/XI8/MM9_g
+ N_VSS_XDFF_Timing_control/XI8/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI8/MM7 N_NOTUSED8_XDFF_Timing_control/XI8/MM7_d
+ N_XDFF_TIMING_CONTROL/XI8/NET71_XDFF_Timing_control/XI8/MM7_g
+ N_VSS_XDFF_Timing_control/XI8/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI8/MM1
+ N_XDFF_TIMING_CONTROL/XI8/NET92_XDFF_Timing_control/XI8/MM1_d
+ N_A<8>_XDFF_Timing_control/XI8/MM1_g N_VDD_XDFF_Timing_control/XI8/MM1_s
+ N_VDD_XDFF_Timing_control/XI8/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI8/MM12
+ N_XDFF_TIMING_CONTROL/XI8/NET92_XDFF_Timing_control/XI8/MM12_d
+ N_CLK_XDFF_Timing_control/XI8/MM12_g
+ N_XDFF_TIMING_CONTROL/XI8/NET75_XDFF_Timing_control/XI8/MM12_s
+ N_VDD_XDFF_Timing_control/XI8/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI8/MM2
+ N_XDFF_TIMING_CONTROL/XI8/NET22_XDFF_Timing_control/XI8/MM2_d
+ N_XDFF_TIMING_CONTROL/XI8/NET75_XDFF_Timing_control/XI8/MM2_g
+ N_VDD_XDFF_Timing_control/XI8/MM2_s N_VDD_XDFF_Timing_control/XI8/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI8/MM15
+ N_XDFF_TIMING_CONTROL/XI8/NET75_XDFF_Timing_control/XI8/MM15_d
+ N_XDFF_TIMING_CONTROL/XI8/NET22_XDFF_Timing_control/XI8/MM15_g
+ N_XDFF_TIMING_CONTROL/XI8/NET23_XDFF_Timing_control/XI8/MM15_s
+ N_VDD_XDFF_Timing_control/XI8/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI8/MM19
+ N_XDFF_TIMING_CONTROL/XI8/NET23_XDFF_Timing_control/XI8/MM19_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI8/MM19_g
+ N_VDD_XDFF_Timing_control/XI8/MM19_s N_VDD_XDFF_Timing_control/XI8/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI8/MM11
+ N_XDFF_TIMING_CONTROL/XI8/NET22_XDFF_Timing_control/XI8/MM11_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI8/MM11_g
+ N_XDFF_TIMING_CONTROL/XI8/NET71_XDFF_Timing_control/XI8/MM11_s
+ N_VDD_XDFF_Timing_control/XI8/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI8/MM5
+ N_XDFF_TIMING_CONTROL/XI8/NET10_XDFF_Timing_control/XI8/MM5_d
+ N_XDFF_TIMING_CONTROL/XI8/NET71_XDFF_Timing_control/XI8/MM5_g
+ N_VDD_XDFF_Timing_control/XI8/MM5_s N_VDD_XDFF_Timing_control/XI8/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI8/MM23
+ N_XDFF_TIMING_CONTROL/XI8/NET71_XDFF_Timing_control/XI8/MM23_d
+ N_XDFF_TIMING_CONTROL/XI8/NET10_XDFF_Timing_control/XI8/MM23_g
+ N_XDFF_TIMING_CONTROL/XI8/NET12_XDFF_Timing_control/XI8/MM23_s
+ N_VDD_XDFF_Timing_control/XI8/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI8/MM22
+ N_XDFF_TIMING_CONTROL/XI8/NET12_XDFF_Timing_control/XI8/MM22_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI8/MM22_g
+ N_VDD_XDFF_Timing_control/XI8/MM22_s N_VDD_XDFF_Timing_control/XI8/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI8/MM8 N_Y_SEL_FF<2>_XDFF_Timing_control/XI8/MM8_d
+ N_XDFF_TIMING_CONTROL/XI8/NET10_XDFF_Timing_control/XI8/MM8_g
+ N_VDD_XDFF_Timing_control/XI8/MM8_s N_VDD_XDFF_Timing_control/XI8/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI8/MM6 N_NOTUSED8_XDFF_Timing_control/XI8/MM6_d
+ N_XDFF_TIMING_CONTROL/XI8/NET71_XDFF_Timing_control/XI8/MM6_g
+ N_VDD_XDFF_Timing_control/XI8/MM6_s N_VDD_XDFF_Timing_control/XI8/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI2/MM0
+ N_XDFF_TIMING_CONTROL/XI2/NET92_XDFF_Timing_control/XI2/MM0_d
+ N_A<1>_XDFF_Timing_control/XI2/MM0_g N_VSS_XDFF_Timing_control/XI2/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI2/MM10
+ N_XDFF_TIMING_CONTROL/XI2/NET92_XDFF_Timing_control/XI2/MM10_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI2/MM10_g
+ N_XDFF_TIMING_CONTROL/XI2/NET75_XDFF_Timing_control/XI2/MM10_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI2/MM3
+ N_XDFF_TIMING_CONTROL/XI2/NET22_XDFF_Timing_control/XI2/MM3_d
+ N_XDFF_TIMING_CONTROL/XI2/NET75_XDFF_Timing_control/XI2/MM3_g
+ N_VSS_XDFF_Timing_control/XI2/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI2/MM16
+ N_XDFF_TIMING_CONTROL/XI2/NET75_XDFF_Timing_control/XI2/MM16_d
+ N_XDFF_TIMING_CONTROL/XI2/NET22_XDFF_Timing_control/XI2/MM16_g
+ N_XDFF_TIMING_CONTROL/XI2/NET60_XDFF_Timing_control/XI2/MM16_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI2/MM20
+ N_XDFF_TIMING_CONTROL/XI2/NET60_XDFF_Timing_control/XI2/MM20_d
+ N_CLK_XDFF_Timing_control/XI2/MM20_g N_VSS_XDFF_Timing_control/XI2/MM20_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI2/MM13
+ N_XDFF_TIMING_CONTROL/XI2/NET22_XDFF_Timing_control/XI2/MM13_d
+ N_CLK_XDFF_Timing_control/XI2/MM13_g
+ N_XDFF_TIMING_CONTROL/XI2/NET71_XDFF_Timing_control/XI2/MM13_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI2/MM4
+ N_XDFF_TIMING_CONTROL/XI2/NET10_XDFF_Timing_control/XI2/MM4_d
+ N_XDFF_TIMING_CONTROL/XI2/NET71_XDFF_Timing_control/XI2/MM4_g
+ N_VSS_XDFF_Timing_control/XI2/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI2/MM24
+ N_XDFF_TIMING_CONTROL/XI2/NET71_XDFF_Timing_control/XI2/MM24_d
+ N_XDFF_TIMING_CONTROL/XI2/NET10_XDFF_Timing_control/XI2/MM24_g
+ N_XDFF_TIMING_CONTROL/XI2/NET56_XDFF_Timing_control/XI2/MM24_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI2/MM21
+ N_XDFF_TIMING_CONTROL/XI2/NET56_XDFF_Timing_control/XI2/MM21_d
+ N_CLK_XDFF_Timing_control/XI2/MM21_g N_VSS_XDFF_Timing_control/XI2/MM21_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI2/MM9 N_X_SEL_FF<1>_XDFF_Timing_control/XI2/MM9_d
+ N_XDFF_TIMING_CONTROL/XI2/NET10_XDFF_Timing_control/XI2/MM9_g
+ N_VSS_XDFF_Timing_control/XI2/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI2/MM7 N_NOTUSED1_XDFF_Timing_control/XI2/MM7_d
+ N_XDFF_TIMING_CONTROL/XI2/NET71_XDFF_Timing_control/XI2/MM7_g
+ N_VSS_XDFF_Timing_control/XI2/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI2/MM1
+ N_XDFF_TIMING_CONTROL/XI2/NET92_XDFF_Timing_control/XI2/MM1_d
+ N_A<1>_XDFF_Timing_control/XI2/MM1_g N_VDD_XDFF_Timing_control/XI2/MM1_s
+ N_VDD_XDFF_Timing_control/XI2/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI2/MM12
+ N_XDFF_TIMING_CONTROL/XI2/NET92_XDFF_Timing_control/XI2/MM12_d
+ N_CLK_XDFF_Timing_control/XI2/MM12_g
+ N_XDFF_TIMING_CONTROL/XI2/NET75_XDFF_Timing_control/XI2/MM12_s
+ N_VDD_XDFF_Timing_control/XI2/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI2/MM2
+ N_XDFF_TIMING_CONTROL/XI2/NET22_XDFF_Timing_control/XI2/MM2_d
+ N_XDFF_TIMING_CONTROL/XI2/NET75_XDFF_Timing_control/XI2/MM2_g
+ N_VDD_XDFF_Timing_control/XI2/MM2_s N_VDD_XDFF_Timing_control/XI2/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI2/MM15
+ N_XDFF_TIMING_CONTROL/XI2/NET75_XDFF_Timing_control/XI2/MM15_d
+ N_XDFF_TIMING_CONTROL/XI2/NET22_XDFF_Timing_control/XI2/MM15_g
+ N_XDFF_TIMING_CONTROL/XI2/NET23_XDFF_Timing_control/XI2/MM15_s
+ N_VDD_XDFF_Timing_control/XI2/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI2/MM19
+ N_XDFF_TIMING_CONTROL/XI2/NET23_XDFF_Timing_control/XI2/MM19_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI2/MM19_g
+ N_VDD_XDFF_Timing_control/XI2/MM19_s N_VDD_XDFF_Timing_control/XI2/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI2/MM11
+ N_XDFF_TIMING_CONTROL/XI2/NET22_XDFF_Timing_control/XI2/MM11_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI2/MM11_g
+ N_XDFF_TIMING_CONTROL/XI2/NET71_XDFF_Timing_control/XI2/MM11_s
+ N_VDD_XDFF_Timing_control/XI2/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI2/MM5
+ N_XDFF_TIMING_CONTROL/XI2/NET10_XDFF_Timing_control/XI2/MM5_d
+ N_XDFF_TIMING_CONTROL/XI2/NET71_XDFF_Timing_control/XI2/MM5_g
+ N_VDD_XDFF_Timing_control/XI2/MM5_s N_VDD_XDFF_Timing_control/XI2/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI2/MM23
+ N_XDFF_TIMING_CONTROL/XI2/NET71_XDFF_Timing_control/XI2/MM23_d
+ N_XDFF_TIMING_CONTROL/XI2/NET10_XDFF_Timing_control/XI2/MM23_g
+ N_XDFF_TIMING_CONTROL/XI2/NET12_XDFF_Timing_control/XI2/MM23_s
+ N_VDD_XDFF_Timing_control/XI2/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI2/MM22
+ N_XDFF_TIMING_CONTROL/XI2/NET12_XDFF_Timing_control/XI2/MM22_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI2/MM22_g
+ N_VDD_XDFF_Timing_control/XI2/MM22_s N_VDD_XDFF_Timing_control/XI2/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI2/MM8 N_X_SEL_FF<1>_XDFF_Timing_control/XI2/MM8_d
+ N_XDFF_TIMING_CONTROL/XI2/NET10_XDFF_Timing_control/XI2/MM8_g
+ N_VDD_XDFF_Timing_control/XI2/MM8_s N_VDD_XDFF_Timing_control/XI2/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI2/MM6 N_NOTUSED1_XDFF_Timing_control/XI2/MM6_d
+ N_XDFF_TIMING_CONTROL/XI2/NET71_XDFF_Timing_control/XI2/MM6_g
+ N_VDD_XDFF_Timing_control/XI2/MM6_s N_VDD_XDFF_Timing_control/XI2/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI7/MM0
+ N_XDFF_TIMING_CONTROL/XI7/NET92_XDFF_Timing_control/XI7/MM0_d
+ N_A<0>_XDFF_Timing_control/XI7/MM0_g N_VSS_XDFF_Timing_control/XI7/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI7/MM10
+ N_XDFF_TIMING_CONTROL/XI7/NET92_XDFF_Timing_control/XI7/MM10_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI7/MM10_g
+ N_XDFF_TIMING_CONTROL/XI7/NET75_XDFF_Timing_control/XI7/MM10_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI7/MM3
+ N_XDFF_TIMING_CONTROL/XI7/NET22_XDFF_Timing_control/XI7/MM3_d
+ N_XDFF_TIMING_CONTROL/XI7/NET75_XDFF_Timing_control/XI7/MM3_g
+ N_VSS_XDFF_Timing_control/XI7/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI7/MM16
+ N_XDFF_TIMING_CONTROL/XI7/NET75_XDFF_Timing_control/XI7/MM16_d
+ N_XDFF_TIMING_CONTROL/XI7/NET22_XDFF_Timing_control/XI7/MM16_g
+ N_XDFF_TIMING_CONTROL/XI7/NET60_XDFF_Timing_control/XI7/MM16_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI7/MM20
+ N_XDFF_TIMING_CONTROL/XI7/NET60_XDFF_Timing_control/XI7/MM20_d
+ N_CLK_XDFF_Timing_control/XI7/MM20_g N_VSS_XDFF_Timing_control/XI7/MM20_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI7/MM13
+ N_XDFF_TIMING_CONTROL/XI7/NET22_XDFF_Timing_control/XI7/MM13_d
+ N_CLK_XDFF_Timing_control/XI7/MM13_g
+ N_XDFF_TIMING_CONTROL/XI7/NET71_XDFF_Timing_control/XI7/MM13_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI7/MM4
+ N_XDFF_TIMING_CONTROL/XI7/NET10_XDFF_Timing_control/XI7/MM4_d
+ N_XDFF_TIMING_CONTROL/XI7/NET71_XDFF_Timing_control/XI7/MM4_g
+ N_VSS_XDFF_Timing_control/XI7/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI7/MM24
+ N_XDFF_TIMING_CONTROL/XI7/NET71_XDFF_Timing_control/XI7/MM24_d
+ N_XDFF_TIMING_CONTROL/XI7/NET10_XDFF_Timing_control/XI7/MM24_g
+ N_XDFF_TIMING_CONTROL/XI7/NET56_XDFF_Timing_control/XI7/MM24_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI7/MM21
+ N_XDFF_TIMING_CONTROL/XI7/NET56_XDFF_Timing_control/XI7/MM21_d
+ N_CLK_XDFF_Timing_control/XI7/MM21_g N_VSS_XDFF_Timing_control/XI7/MM21_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI7/MM9 N_X_SEL_FF<0>_XDFF_Timing_control/XI7/MM9_d
+ N_XDFF_TIMING_CONTROL/XI7/NET10_XDFF_Timing_control/XI7/MM9_g
+ N_VSS_XDFF_Timing_control/XI7/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI7/MM7 N_NOTUSED0_XDFF_Timing_control/XI7/MM7_d
+ N_XDFF_TIMING_CONTROL/XI7/NET71_XDFF_Timing_control/XI7/MM7_g
+ N_VSS_XDFF_Timing_control/XI7/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI7/MM1
+ N_XDFF_TIMING_CONTROL/XI7/NET92_XDFF_Timing_control/XI7/MM1_d
+ N_A<0>_XDFF_Timing_control/XI7/MM1_g N_VDD_XDFF_Timing_control/XI7/MM1_s
+ N_VDD_XDFF_Timing_control/XI7/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI7/MM12
+ N_XDFF_TIMING_CONTROL/XI7/NET92_XDFF_Timing_control/XI7/MM12_d
+ N_CLK_XDFF_Timing_control/XI7/MM12_g
+ N_XDFF_TIMING_CONTROL/XI7/NET75_XDFF_Timing_control/XI7/MM12_s
+ N_VDD_XDFF_Timing_control/XI7/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI7/MM2
+ N_XDFF_TIMING_CONTROL/XI7/NET22_XDFF_Timing_control/XI7/MM2_d
+ N_XDFF_TIMING_CONTROL/XI7/NET75_XDFF_Timing_control/XI7/MM2_g
+ N_VDD_XDFF_Timing_control/XI7/MM2_s N_VDD_XDFF_Timing_control/XI7/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI7/MM15
+ N_XDFF_TIMING_CONTROL/XI7/NET75_XDFF_Timing_control/XI7/MM15_d
+ N_XDFF_TIMING_CONTROL/XI7/NET22_XDFF_Timing_control/XI7/MM15_g
+ N_XDFF_TIMING_CONTROL/XI7/NET23_XDFF_Timing_control/XI7/MM15_s
+ N_VDD_XDFF_Timing_control/XI7/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI7/MM19
+ N_XDFF_TIMING_CONTROL/XI7/NET23_XDFF_Timing_control/XI7/MM19_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI7/MM19_g
+ N_VDD_XDFF_Timing_control/XI7/MM19_s N_VDD_XDFF_Timing_control/XI7/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI7/MM11
+ N_XDFF_TIMING_CONTROL/XI7/NET22_XDFF_Timing_control/XI7/MM11_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI7/MM11_g
+ N_XDFF_TIMING_CONTROL/XI7/NET71_XDFF_Timing_control/XI7/MM11_s
+ N_VDD_XDFF_Timing_control/XI7/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI7/MM5
+ N_XDFF_TIMING_CONTROL/XI7/NET10_XDFF_Timing_control/XI7/MM5_d
+ N_XDFF_TIMING_CONTROL/XI7/NET71_XDFF_Timing_control/XI7/MM5_g
+ N_VDD_XDFF_Timing_control/XI7/MM5_s N_VDD_XDFF_Timing_control/XI7/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI7/MM23
+ N_XDFF_TIMING_CONTROL/XI7/NET71_XDFF_Timing_control/XI7/MM23_d
+ N_XDFF_TIMING_CONTROL/XI7/NET10_XDFF_Timing_control/XI7/MM23_g
+ N_XDFF_TIMING_CONTROL/XI7/NET12_XDFF_Timing_control/XI7/MM23_s
+ N_VDD_XDFF_Timing_control/XI7/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI7/MM22
+ N_XDFF_TIMING_CONTROL/XI7/NET12_XDFF_Timing_control/XI7/MM22_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI7/MM22_g
+ N_VDD_XDFF_Timing_control/XI7/MM22_s N_VDD_XDFF_Timing_control/XI7/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI7/MM8 N_X_SEL_FF<0>_XDFF_Timing_control/XI7/MM8_d
+ N_XDFF_TIMING_CONTROL/XI7/NET10_XDFF_Timing_control/XI7/MM8_g
+ N_VDD_XDFF_Timing_control/XI7/MM8_s N_VDD_XDFF_Timing_control/XI7/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI7/MM6 N_NOTUSED0_XDFF_Timing_control/XI7/MM6_d
+ N_XDFF_TIMING_CONTROL/XI7/NET71_XDFF_Timing_control/XI7/MM6_g
+ N_VDD_XDFF_Timing_control/XI7/MM6_s N_VDD_XDFF_Timing_control/XI7/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI4/MM0
+ N_XDFF_TIMING_CONTROL/XI4/NET92_XDFF_Timing_control/XI4/MM0_d
+ N_A<3>_XDFF_Timing_control/XI4/MM0_g N_VSS_XDFF_Timing_control/XI4/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI4/MM10
+ N_XDFF_TIMING_CONTROL/XI4/NET92_XDFF_Timing_control/XI4/MM10_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI4/MM10_g
+ N_XDFF_TIMING_CONTROL/XI4/NET75_XDFF_Timing_control/XI4/MM10_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI4/MM3
+ N_XDFF_TIMING_CONTROL/XI4/NET22_XDFF_Timing_control/XI4/MM3_d
+ N_XDFF_TIMING_CONTROL/XI4/NET75_XDFF_Timing_control/XI4/MM3_g
+ N_VSS_XDFF_Timing_control/XI4/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI4/MM16
+ N_XDFF_TIMING_CONTROL/XI4/NET75_XDFF_Timing_control/XI4/MM16_d
+ N_XDFF_TIMING_CONTROL/XI4/NET22_XDFF_Timing_control/XI4/MM16_g
+ N_XDFF_TIMING_CONTROL/XI4/NET60_XDFF_Timing_control/XI4/MM16_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI4/MM20
+ N_XDFF_TIMING_CONTROL/XI4/NET60_XDFF_Timing_control/XI4/MM20_d
+ N_CLK_XDFF_Timing_control/XI4/MM20_g N_VSS_XDFF_Timing_control/XI4/MM20_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI4/MM13
+ N_XDFF_TIMING_CONTROL/XI4/NET22_XDFF_Timing_control/XI4/MM13_d
+ N_CLK_XDFF_Timing_control/XI4/MM13_g
+ N_XDFF_TIMING_CONTROL/XI4/NET71_XDFF_Timing_control/XI4/MM13_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI4/MM4
+ N_XDFF_TIMING_CONTROL/XI4/NET10_XDFF_Timing_control/XI4/MM4_d
+ N_XDFF_TIMING_CONTROL/XI4/NET71_XDFF_Timing_control/XI4/MM4_g
+ N_VSS_XDFF_Timing_control/XI4/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI4/MM24
+ N_XDFF_TIMING_CONTROL/XI4/NET71_XDFF_Timing_control/XI4/MM24_d
+ N_XDFF_TIMING_CONTROL/XI4/NET10_XDFF_Timing_control/XI4/MM24_g
+ N_XDFF_TIMING_CONTROL/XI4/NET56_XDFF_Timing_control/XI4/MM24_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI4/MM21
+ N_XDFF_TIMING_CONTROL/XI4/NET56_XDFF_Timing_control/XI4/MM21_d
+ N_CLK_XDFF_Timing_control/XI4/MM21_g N_VSS_XDFF_Timing_control/XI4/MM21_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI4/MM9 N_X_SEL_FF<3>_XDFF_Timing_control/XI4/MM9_d
+ N_XDFF_TIMING_CONTROL/XI4/NET10_XDFF_Timing_control/XI4/MM9_g
+ N_VSS_XDFF_Timing_control/XI4/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI4/MM7 N_NOTUSED3_XDFF_Timing_control/XI4/MM7_d
+ N_XDFF_TIMING_CONTROL/XI4/NET71_XDFF_Timing_control/XI4/MM7_g
+ N_VSS_XDFF_Timing_control/XI4/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI4/MM1
+ N_XDFF_TIMING_CONTROL/XI4/NET92_XDFF_Timing_control/XI4/MM1_d
+ N_A<3>_XDFF_Timing_control/XI4/MM1_g N_VDD_XDFF_Timing_control/XI4/MM1_s
+ N_VDD_XDFF_Timing_control/XI4/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI4/MM12
+ N_XDFF_TIMING_CONTROL/XI4/NET92_XDFF_Timing_control/XI4/MM12_d
+ N_CLK_XDFF_Timing_control/XI4/MM12_g
+ N_XDFF_TIMING_CONTROL/XI4/NET75_XDFF_Timing_control/XI4/MM12_s
+ N_VDD_XDFF_Timing_control/XI4/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI4/MM2
+ N_XDFF_TIMING_CONTROL/XI4/NET22_XDFF_Timing_control/XI4/MM2_d
+ N_XDFF_TIMING_CONTROL/XI4/NET75_XDFF_Timing_control/XI4/MM2_g
+ N_VDD_XDFF_Timing_control/XI4/MM2_s N_VDD_XDFF_Timing_control/XI4/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI4/MM15
+ N_XDFF_TIMING_CONTROL/XI4/NET75_XDFF_Timing_control/XI4/MM15_d
+ N_XDFF_TIMING_CONTROL/XI4/NET22_XDFF_Timing_control/XI4/MM15_g
+ N_XDFF_TIMING_CONTROL/XI4/NET23_XDFF_Timing_control/XI4/MM15_s
+ N_VDD_XDFF_Timing_control/XI4/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI4/MM19
+ N_XDFF_TIMING_CONTROL/XI4/NET23_XDFF_Timing_control/XI4/MM19_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI4/MM19_g
+ N_VDD_XDFF_Timing_control/XI4/MM19_s N_VDD_XDFF_Timing_control/XI4/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI4/MM11
+ N_XDFF_TIMING_CONTROL/XI4/NET22_XDFF_Timing_control/XI4/MM11_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI4/MM11_g
+ N_XDFF_TIMING_CONTROL/XI4/NET71_XDFF_Timing_control/XI4/MM11_s
+ N_VDD_XDFF_Timing_control/XI4/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI4/MM5
+ N_XDFF_TIMING_CONTROL/XI4/NET10_XDFF_Timing_control/XI4/MM5_d
+ N_XDFF_TIMING_CONTROL/XI4/NET71_XDFF_Timing_control/XI4/MM5_g
+ N_VDD_XDFF_Timing_control/XI4/MM5_s N_VDD_XDFF_Timing_control/XI4/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI4/MM23
+ N_XDFF_TIMING_CONTROL/XI4/NET71_XDFF_Timing_control/XI4/MM23_d
+ N_XDFF_TIMING_CONTROL/XI4/NET10_XDFF_Timing_control/XI4/MM23_g
+ N_XDFF_TIMING_CONTROL/XI4/NET12_XDFF_Timing_control/XI4/MM23_s
+ N_VDD_XDFF_Timing_control/XI4/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI4/MM22
+ N_XDFF_TIMING_CONTROL/XI4/NET12_XDFF_Timing_control/XI4/MM22_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI4/MM22_g
+ N_VDD_XDFF_Timing_control/XI4/MM22_s N_VDD_XDFF_Timing_control/XI4/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI4/MM8 N_X_SEL_FF<3>_XDFF_Timing_control/XI4/MM8_d
+ N_XDFF_TIMING_CONTROL/XI4/NET10_XDFF_Timing_control/XI4/MM8_g
+ N_VDD_XDFF_Timing_control/XI4/MM8_s N_VDD_XDFF_Timing_control/XI4/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI4/MM6 N_NOTUSED3_XDFF_Timing_control/XI4/MM6_d
+ N_XDFF_TIMING_CONTROL/XI4/NET71_XDFF_Timing_control/XI4/MM6_g
+ N_VDD_XDFF_Timing_control/XI4/MM6_s N_VDD_XDFF_Timing_control/XI4/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI5/MM0
+ N_XDFF_TIMING_CONTROL/XI5/NET92_XDFF_Timing_control/XI5/MM0_d
+ N_A<4>_XDFF_Timing_control/XI5/MM0_g N_VSS_XDFF_Timing_control/XI5/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI5/MM10
+ N_XDFF_TIMING_CONTROL/XI5/NET92_XDFF_Timing_control/XI5/MM10_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI5/MM10_g
+ N_XDFF_TIMING_CONTROL/XI5/NET75_XDFF_Timing_control/XI5/MM10_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI5/MM3
+ N_XDFF_TIMING_CONTROL/XI5/NET22_XDFF_Timing_control/XI5/MM3_d
+ N_XDFF_TIMING_CONTROL/XI5/NET75_XDFF_Timing_control/XI5/MM3_g
+ N_VSS_XDFF_Timing_control/XI5/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI5/MM16
+ N_XDFF_TIMING_CONTROL/XI5/NET75_XDFF_Timing_control/XI5/MM16_d
+ N_XDFF_TIMING_CONTROL/XI5/NET22_XDFF_Timing_control/XI5/MM16_g
+ N_XDFF_TIMING_CONTROL/XI5/NET60_XDFF_Timing_control/XI5/MM16_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI5/MM20
+ N_XDFF_TIMING_CONTROL/XI5/NET60_XDFF_Timing_control/XI5/MM20_d
+ N_CLK_XDFF_Timing_control/XI5/MM20_g N_VSS_XDFF_Timing_control/XI5/MM20_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI5/MM13
+ N_XDFF_TIMING_CONTROL/XI5/NET22_XDFF_Timing_control/XI5/MM13_d
+ N_CLK_XDFF_Timing_control/XI5/MM13_g
+ N_XDFF_TIMING_CONTROL/XI5/NET71_XDFF_Timing_control/XI5/MM13_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXDFF_Timing_control/XI5/MM4
+ N_XDFF_TIMING_CONTROL/XI5/NET10_XDFF_Timing_control/XI5/MM4_d
+ N_XDFF_TIMING_CONTROL/XI5/NET71_XDFF_Timing_control/XI5/MM4_g
+ N_VSS_XDFF_Timing_control/XI5/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI5/MM24
+ N_XDFF_TIMING_CONTROL/XI5/NET71_XDFF_Timing_control/XI5/MM24_d
+ N_XDFF_TIMING_CONTROL/XI5/NET10_XDFF_Timing_control/XI5/MM24_g
+ N_XDFF_TIMING_CONTROL/XI5/NET56_XDFF_Timing_control/XI5/MM24_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI5/MM21
+ N_XDFF_TIMING_CONTROL/XI5/NET56_XDFF_Timing_control/XI5/MM21_d
+ N_CLK_XDFF_Timing_control/XI5/MM21_g N_VSS_XDFF_Timing_control/XI5/MM21_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI5/MM9 N_X_SEL_FF<4>_XDFF_Timing_control/XI5/MM9_d
+ N_XDFF_TIMING_CONTROL/XI5/NET10_XDFF_Timing_control/XI5/MM9_g
+ N_VSS_XDFF_Timing_control/XI5/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI5/MM7 N_NOTUSED4_XDFF_Timing_control/XI5/MM7_d
+ N_XDFF_TIMING_CONTROL/XI5/NET71_XDFF_Timing_control/XI5/MM7_g
+ N_VSS_XDFF_Timing_control/XI5/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXDFF_Timing_control/XI5/MM1
+ N_XDFF_TIMING_CONTROL/XI5/NET92_XDFF_Timing_control/XI5/MM1_d
+ N_A<4>_XDFF_Timing_control/XI5/MM1_g N_VDD_XDFF_Timing_control/XI5/MM1_s
+ N_VDD_XDFF_Timing_control/XI5/MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI5/MM12
+ N_XDFF_TIMING_CONTROL/XI5/NET92_XDFF_Timing_control/XI5/MM12_d
+ N_CLK_XDFF_Timing_control/XI5/MM12_g
+ N_XDFF_TIMING_CONTROL/XI5/NET75_XDFF_Timing_control/XI5/MM12_s
+ N_VDD_XDFF_Timing_control/XI5/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI5/MM2
+ N_XDFF_TIMING_CONTROL/XI5/NET22_XDFF_Timing_control/XI5/MM2_d
+ N_XDFF_TIMING_CONTROL/XI5/NET75_XDFF_Timing_control/XI5/MM2_g
+ N_VDD_XDFF_Timing_control/XI5/MM2_s N_VDD_XDFF_Timing_control/XI5/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI5/MM15
+ N_XDFF_TIMING_CONTROL/XI5/NET75_XDFF_Timing_control/XI5/MM15_d
+ N_XDFF_TIMING_CONTROL/XI5/NET22_XDFF_Timing_control/XI5/MM15_g
+ N_XDFF_TIMING_CONTROL/XI5/NET23_XDFF_Timing_control/XI5/MM15_s
+ N_VDD_XDFF_Timing_control/XI5/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI5/MM19
+ N_XDFF_TIMING_CONTROL/XI5/NET23_XDFF_Timing_control/XI5/MM19_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI5/MM19_g
+ N_VDD_XDFF_Timing_control/XI5/MM19_s N_VDD_XDFF_Timing_control/XI5/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI5/MM11
+ N_XDFF_TIMING_CONTROL/XI5/NET22_XDFF_Timing_control/XI5/MM11_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI5/MM11_g
+ N_XDFF_TIMING_CONTROL/XI5/NET71_XDFF_Timing_control/XI5/MM11_s
+ N_VDD_XDFF_Timing_control/XI5/MM1_b P_18 L=1.8e-07 W=1e-06 AD=4.9e-13
+ AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXDFF_Timing_control/XI5/MM5
+ N_XDFF_TIMING_CONTROL/XI5/NET10_XDFF_Timing_control/XI5/MM5_d
+ N_XDFF_TIMING_CONTROL/XI5/NET71_XDFF_Timing_control/XI5/MM5_g
+ N_VDD_XDFF_Timing_control/XI5/MM5_s N_VDD_XDFF_Timing_control/XI5/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI5/MM23
+ N_XDFF_TIMING_CONTROL/XI5/NET71_XDFF_Timing_control/XI5/MM23_d
+ N_XDFF_TIMING_CONTROL/XI5/NET10_XDFF_Timing_control/XI5/MM23_g
+ N_XDFF_TIMING_CONTROL/XI5/NET12_XDFF_Timing_control/XI5/MM23_s
+ N_VDD_XDFF_Timing_control/XI5/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXDFF_Timing_control/XI5/MM22
+ N_XDFF_TIMING_CONTROL/XI5/NET12_XDFF_Timing_control/XI5/MM22_d
+ N_XDFF_TIMING_CONTROL/NET28_XDFF_Timing_control/XI5/MM22_g
+ N_VDD_XDFF_Timing_control/XI5/MM22_s N_VDD_XDFF_Timing_control/XI5/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXDFF_Timing_control/XI5/MM8 N_X_SEL_FF<4>_XDFF_Timing_control/XI5/MM8_d
+ N_XDFF_TIMING_CONTROL/XI5/NET10_XDFF_Timing_control/XI5/MM8_g
+ N_VDD_XDFF_Timing_control/XI5/MM8_s N_VDD_XDFF_Timing_control/XI5/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXDFF_Timing_control/XI5/MM6 N_NOTUSED4_XDFF_Timing_control/XI5/MM6_d
+ N_XDFF_TIMING_CONTROL/XI5/NET71_XDFF_Timing_control/XI5/MM6_g
+ N_VDD_XDFF_Timing_control/XI5/MM6_s N_VDD_XDFF_Timing_control/XI5/MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXXDec/XI40/XI17/MN N_XXDEC/XI40/NET22_XXDec/XI40/XI17/MN_d
+ N_X_SEL_FF<0>_XXDec/XI40/XI17/MN_g N_VSS_XXDec/XI40/XI17/MN_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXXDec/XI39/XI17/MN N_XXDEC/XI39/NET22_XXDec/XI39/XI17/MN_d
+ N_X_SEL_FF<3>_XXDec/XI39/XI17/MN_g N_VSS_XXDec/XI39/XI17/MN_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXXDec/XI40/XI18/MN N_XXDEC/XI40/NET18_XXDec/XI40/XI18/MN_d
+ N_X_SEL_FF<1>_XXDec/XI40/XI18/MN_g N_VSS_XXDec/XI40/XI18/MN_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXXDec/XI39/XI18/MN N_XXDEC/XI39/NET18_XXDec/XI39/XI18/MN_d
+ N_X_SEL_FF<4>_XXDec/XI39/XI18/MN_g N_VSS_XXDec/XI39/XI18/MN_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXXDec/XI40/XI19/MN N_XXDEC/XI40/NET14_XXDec/XI40/XI19/MN_d
+ N_X_SEL_FF<2>_XXDec/XI40/XI19/MN_g N_VSS_XXDec/XI40/XI19/MN_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXXDec/XI39/XI19/MN N_XXDEC/XI39/NET14_XXDec/XI39/XI19/MN_d
+ N_X_SEL_FF<5>_XXDec/XI39/XI19/MN_g N_VSS_XXDec/XI39/XI19/MN_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXXDec/XI40/XI26/MM3 N_XXDEC/XI40/XI26/NET24_XXDec/XI40/XI26/MM3_d
+ N_WL_EN_XXDec/XI40/XI26/MM3_g N_VSS_XXDec/XI40/XI26/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI40/XI25/MM3 N_XXDEC/XI40/XI25/NET24_XXDec/XI40/XI25/MM3_d
+ N_WL_EN_XXDec/XI40/XI25/MM3_g N_VSS_XXDec/XI40/XI25/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI40/XI22/MM3 N_XXDEC/XI40/XI22/NET24_XXDec/XI40/XI22/MM3_d
+ N_WL_EN_XXDec/XI40/XI22/MM3_g N_VSS_XXDec/XI40/XI22/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI40/XI21/MM3 N_XXDEC/XI40/XI21/NET24_XXDec/XI40/XI21/MM3_d
+ N_WL_EN_XXDec/XI40/XI21/MM3_g N_VSS_XXDec/XI40/XI21/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI39/XI21/MM3 N_XXDEC/XI39/XI21/NET24_XXDec/XI39/XI21/MM3_d
+ N_WL_EN_XXDec/XI39/XI21/MM3_g N_VSS_XXDec/XI39/XI21/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI39/XI22/MM3 N_XXDEC/XI39/XI22/NET24_XXDec/XI39/XI22/MM3_d
+ N_WL_EN_XXDec/XI39/XI22/MM3_g N_VSS_XXDec/XI39/XI22/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI39/XI25/MM3 N_XXDEC/XI39/XI25/NET24_XXDec/XI39/XI25/MM3_d
+ N_WL_EN_XXDec/XI39/XI25/MM3_g N_VSS_XXDec/XI39/XI25/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI39/XI26/MM3 N_XXDEC/XI39/XI26/NET24_XXDec/XI39/XI26/MM3_d
+ N_WL_EN_XXDec/XI39/XI26/MM3_g N_VSS_XXDec/XI39/XI26/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI40/XI26/MM2 N_XXDEC/XI40/XI26/NET28_XXDec/XI40/XI26/MM2_d
+ N_XXDEC/XI40/NET14_XXDec/XI40/XI26/MM2_g
+ N_XXDEC/XI40/XI26/NET24_XXDec/XI40/XI26/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI25/MM2 N_XXDEC/XI40/XI25/NET28_XXDec/XI40/XI25/MM2_d
+ N_XXDEC/XI40/NET14_XXDec/XI40/XI25/MM2_g
+ N_XXDEC/XI40/XI25/NET24_XXDec/XI40/XI25/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI22/MM2 N_XXDEC/XI40/XI22/NET28_XXDec/XI40/XI22/MM2_d
+ N_X_SEL_FF<2>_XXDec/XI40/XI22/MM2_g
+ N_XXDEC/XI40/XI22/NET24_XXDec/XI40/XI22/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI21/MM2 N_XXDEC/XI40/XI21/NET28_XXDec/XI40/XI21/MM2_d
+ N_X_SEL_FF<2>_XXDec/XI40/XI21/MM2_g
+ N_XXDEC/XI40/XI21/NET24_XXDec/XI40/XI21/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI21/MM2 N_XXDEC/XI39/XI21/NET28_XXDec/XI39/XI21/MM2_d
+ N_X_SEL_FF<5>_XXDec/XI39/XI21/MM2_g
+ N_XXDEC/XI39/XI21/NET24_XXDec/XI39/XI21/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI22/MM2 N_XXDEC/XI39/XI22/NET28_XXDec/XI39/XI22/MM2_d
+ N_X_SEL_FF<5>_XXDec/XI39/XI22/MM2_g
+ N_XXDEC/XI39/XI22/NET24_XXDec/XI39/XI22/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI25/MM2 N_XXDEC/XI39/XI25/NET28_XXDec/XI39/XI25/MM2_d
+ N_XXDEC/XI39/NET14_XXDec/XI39/XI25/MM2_g
+ N_XXDEC/XI39/XI25/NET24_XXDec/XI39/XI25/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI26/MM2 N_XXDEC/XI39/XI26/NET28_XXDec/XI39/XI26/MM2_d
+ N_XXDEC/XI39/NET14_XXDec/XI39/XI26/MM2_g
+ N_XXDEC/XI39/XI26/NET24_XXDec/XI39/XI26/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI26/MM1 N_XXDEC/XI40/XI26/NET32_XXDec/XI40/XI26/MM1_d
+ N_XXDEC/XI40/NET18_XXDec/XI40/XI26/MM1_g
+ N_XXDEC/XI40/XI26/NET28_XXDec/XI40/XI26/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI25/MM1 N_XXDEC/XI40/XI25/NET32_XXDec/XI40/XI25/MM1_d
+ N_X_SEL_FF<1>_XXDec/XI40/XI25/MM1_g
+ N_XXDEC/XI40/XI25/NET28_XXDec/XI40/XI25/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI22/MM1 N_XXDEC/XI40/XI22/NET32_XXDec/XI40/XI22/MM1_d
+ N_XXDEC/XI40/NET18_XXDec/XI40/XI22/MM1_g
+ N_XXDEC/XI40/XI22/NET28_XXDec/XI40/XI22/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI21/MM1 N_XXDEC/XI40/XI21/NET32_XXDec/XI40/XI21/MM1_d
+ N_X_SEL_FF<1>_XXDec/XI40/XI21/MM1_g
+ N_XXDEC/XI40/XI21/NET28_XXDec/XI40/XI21/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI21/MM1 N_XXDEC/XI39/XI21/NET32_XXDec/XI39/XI21/MM1_d
+ N_X_SEL_FF<4>_XXDec/XI39/XI21/MM1_g
+ N_XXDEC/XI39/XI21/NET28_XXDec/XI39/XI21/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI22/MM1 N_XXDEC/XI39/XI22/NET32_XXDec/XI39/XI22/MM1_d
+ N_XXDEC/XI39/NET18_XXDec/XI39/XI22/MM1_g
+ N_XXDEC/XI39/XI22/NET28_XXDec/XI39/XI22/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI25/MM1 N_XXDEC/XI39/XI25/NET32_XXDec/XI39/XI25/MM1_d
+ N_X_SEL_FF<4>_XXDec/XI39/XI25/MM1_g
+ N_XXDEC/XI39/XI25/NET28_XXDec/XI39/XI25/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI26/MM1 N_XXDEC/XI39/XI26/NET32_XXDec/XI39/XI26/MM1_d
+ N_XXDEC/XI39/NET18_XXDec/XI39/XI26/MM1_g
+ N_XXDEC/XI39/XI26/NET28_XXDec/XI39/XI26/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI26/MM0 N_XXDEC/NET0143_XXDec/XI40/XI26/MM0_d
+ N_X_SEL_FF<0>_XXDec/XI40/XI26/MM0_g
+ N_XXDEC/XI40/XI26/NET32_XXDec/XI40/XI26/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI25/MM0 N_XXDEC/NET0142_XXDec/XI40/XI25/MM0_d
+ N_XXDEC/XI40/NET22_XXDec/XI40/XI25/MM0_g
+ N_XXDEC/XI40/XI25/NET32_XXDec/XI40/XI25/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI22/MM0 N_XXDEC/NET0139_XXDec/XI40/XI22/MM0_d
+ N_X_SEL_FF<0>_XXDec/XI40/XI22/MM0_g
+ N_XXDEC/XI40/XI22/NET32_XXDec/XI40/XI22/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI21/MM0 N_XXDEC/NET0138_XXDec/XI40/XI21/MM0_d
+ N_XXDEC/XI40/NET22_XXDec/XI40/XI21/MM0_g
+ N_XXDEC/XI40/XI21/NET32_XXDec/XI40/XI21/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI21/MM0 N_XXDEC/NET187_XXDec/XI39/XI21/MM0_d
+ N_XXDEC/XI39/NET22_XXDec/XI39/XI21/MM0_g
+ N_XXDEC/XI39/XI21/NET32_XXDec/XI39/XI21/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI22/MM0 N_XXDEC/NET188_XXDec/XI39/XI22/MM0_d
+ N_X_SEL_FF<3>_XXDec/XI39/XI22/MM0_g
+ N_XXDEC/XI39/XI22/NET32_XXDec/XI39/XI22/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI25/MM0 N_XXDEC/NET0220_XXDec/XI39/XI25/MM0_d
+ N_XXDEC/XI39/NET22_XXDec/XI39/XI25/MM0_g
+ N_XXDEC/XI39/XI25/NET32_XXDec/XI39/XI25/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI26/MM0 N_XXDEC/NET192_XXDec/XI39/XI26/MM0_d
+ N_X_SEL_FF<3>_XXDec/XI39/XI26/MM0_g
+ N_XXDEC/XI39/XI26/NET32_XXDec/XI39/XI26/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI27/MM3 N_XXDEC/XI40/XI27/NET24_XXDec/XI40/XI27/MM3_d
+ N_WL_EN_XXDec/XI40/XI27/MM3_g N_VSS_XXDec/XI40/XI27/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI40/XI24/MM3 N_XXDEC/XI40/XI24/NET24_XXDec/XI40/XI24/MM3_d
+ N_WL_EN_XXDec/XI40/XI24/MM3_g N_VSS_XXDec/XI40/XI24/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI40/XI23/MM3 N_XXDEC/XI40/XI23/NET24_XXDec/XI40/XI23/MM3_d
+ N_WL_EN_XXDec/XI40/XI23/MM3_g N_VSS_XXDec/XI40/XI23/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI40/XI20/MM3 N_XXDEC/XI40/XI20/NET24_XXDec/XI40/XI20/MM3_d
+ N_WL_EN_XXDec/XI40/XI20/MM3_g N_VSS_XXDec/XI40/XI20/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI39/XI20/MM3 N_XXDEC/XI39/XI20/NET24_XXDec/XI39/XI20/MM3_d
+ N_WL_EN_XXDec/XI39/XI20/MM3_g N_VSS_XXDec/XI39/XI20/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI39/XI23/MM3 N_XXDEC/XI39/XI23/NET24_XXDec/XI39/XI23/MM3_d
+ N_WL_EN_XXDec/XI39/XI23/MM3_g N_VSS_XXDec/XI39/XI23/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI39/XI24/MM3 N_XXDEC/XI39/XI24/NET24_XXDec/XI39/XI24/MM3_d
+ N_WL_EN_XXDec/XI39/XI24/MM3_g N_VSS_XXDec/XI39/XI24/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI39/XI27/MM3 N_XXDEC/XI39/XI27/NET24_XXDec/XI39/XI27/MM3_d
+ N_WL_EN_XXDec/XI39/XI27/MM3_g N_VSS_XXDec/XI39/XI27/MM3_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=2.45e-13 PD=5.1e-07 PS=1.48e-06
mXXDec/XI40/XI27/MM2 N_XXDEC/XI40/XI27/NET28_XXDec/XI40/XI27/MM2_d
+ N_XXDEC/XI40/NET14_XXDec/XI40/XI27/MM2_g
+ N_XXDEC/XI40/XI27/NET24_XXDec/XI40/XI27/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI24/MM2 N_XXDEC/XI40/XI24/NET28_XXDec/XI40/XI24/MM2_d
+ N_XXDEC/XI40/NET14_XXDec/XI40/XI24/MM2_g
+ N_XXDEC/XI40/XI24/NET24_XXDec/XI40/XI24/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI23/MM2 N_XXDEC/XI40/XI23/NET28_XXDec/XI40/XI23/MM2_d
+ N_X_SEL_FF<2>_XXDec/XI40/XI23/MM2_g
+ N_XXDEC/XI40/XI23/NET24_XXDec/XI40/XI23/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI20/MM2 N_XXDEC/XI40/XI20/NET28_XXDec/XI40/XI20/MM2_d
+ N_X_SEL_FF<2>_XXDec/XI40/XI20/MM2_g
+ N_XXDEC/XI40/XI20/NET24_XXDec/XI40/XI20/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI20/MM2 N_XXDEC/XI39/XI20/NET28_XXDec/XI39/XI20/MM2_d
+ N_X_SEL_FF<5>_XXDec/XI39/XI20/MM2_g
+ N_XXDEC/XI39/XI20/NET24_XXDec/XI39/XI20/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI23/MM2 N_XXDEC/XI39/XI23/NET28_XXDec/XI39/XI23/MM2_d
+ N_X_SEL_FF<5>_XXDec/XI39/XI23/MM2_g
+ N_XXDEC/XI39/XI23/NET24_XXDec/XI39/XI23/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI24/MM2 N_XXDEC/XI39/XI24/NET28_XXDec/XI39/XI24/MM2_d
+ N_XXDEC/XI39/NET14_XXDec/XI39/XI24/MM2_g
+ N_XXDEC/XI39/XI24/NET24_XXDec/XI39/XI24/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI27/MM2 N_XXDEC/XI39/XI27/NET28_XXDec/XI39/XI27/MM2_d
+ N_XXDEC/XI39/NET14_XXDec/XI39/XI27/MM2_g
+ N_XXDEC/XI39/XI27/NET24_XXDec/XI39/XI27/MM2_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI27/MM1 N_XXDEC/XI40/XI27/NET32_XXDec/XI40/XI27/MM1_d
+ N_XXDEC/XI40/NET18_XXDec/XI40/XI27/MM1_g
+ N_XXDEC/XI40/XI27/NET28_XXDec/XI40/XI27/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI24/MM1 N_XXDEC/XI40/XI24/NET32_XXDec/XI40/XI24/MM1_d
+ N_X_SEL_FF<1>_XXDec/XI40/XI24/MM1_g
+ N_XXDEC/XI40/XI24/NET28_XXDec/XI40/XI24/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI23/MM1 N_XXDEC/XI40/XI23/NET32_XXDec/XI40/XI23/MM1_d
+ N_XXDEC/XI40/NET18_XXDec/XI40/XI23/MM1_g
+ N_XXDEC/XI40/XI23/NET28_XXDec/XI40/XI23/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI20/MM1 N_XXDEC/XI40/XI20/NET32_XXDec/XI40/XI20/MM1_d
+ N_X_SEL_FF<1>_XXDec/XI40/XI20/MM1_g
+ N_XXDEC/XI40/XI20/NET28_XXDec/XI40/XI20/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI20/MM1 N_XXDEC/XI39/XI20/NET32_XXDec/XI39/XI20/MM1_d
+ N_X_SEL_FF<4>_XXDec/XI39/XI20/MM1_g
+ N_XXDEC/XI39/XI20/NET28_XXDec/XI39/XI20/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI23/MM1 N_XXDEC/XI39/XI23/NET32_XXDec/XI39/XI23/MM1_d
+ N_XXDEC/XI39/NET18_XXDec/XI39/XI23/MM1_g
+ N_XXDEC/XI39/XI23/NET28_XXDec/XI39/XI23/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI24/MM1 N_XXDEC/XI39/XI24/NET32_XXDec/XI39/XI24/MM1_d
+ N_X_SEL_FF<4>_XXDec/XI39/XI24/MM1_g
+ N_XXDEC/XI39/XI24/NET28_XXDec/XI39/XI24/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI27/MM1 N_XXDEC/XI39/XI27/NET32_XXDec/XI39/XI27/MM1_d
+ N_XXDEC/XI39/NET18_XXDec/XI39/XI27/MM1_g
+ N_XXDEC/XI39/XI27/NET28_XXDec/XI39/XI27/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.275e-13
+ AS=1.275e-13 PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI27/MM0 N_XXDEC/NET0144_XXDec/XI40/XI27/MM0_d
+ N_XXDEC/XI40/NET22_XXDec/XI40/XI27/MM0_g
+ N_XXDEC/XI40/XI27/NET32_XXDec/XI40/XI27/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI24/MM0 N_XXDEC/NET0141_XXDec/XI40/XI24/MM0_d
+ N_X_SEL_FF<0>_XXDec/XI40/XI24/MM0_g
+ N_XXDEC/XI40/XI24/NET32_XXDec/XI40/XI24/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI23/MM0 N_XXDEC/NET0140_XXDec/XI40/XI23/MM0_d
+ N_XXDEC/XI40/NET22_XXDec/XI40/XI23/MM0_g
+ N_XXDEC/XI40/XI23/NET32_XXDec/XI40/XI23/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI20/MM0 N_XXDEC/NET0137_XXDec/XI40/XI20/MM0_d
+ N_X_SEL_FF<0>_XXDec/XI40/XI20/MM0_g
+ N_XXDEC/XI40/XI20/NET32_XXDec/XI40/XI20/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI20/MM0 N_XXDEC/NET0123_XXDec/XI39/XI20/MM0_d
+ N_X_SEL_FF<3>_XXDec/XI39/XI20/MM0_g
+ N_XXDEC/XI39/XI20/NET32_XXDec/XI39/XI20/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI23/MM0 N_XXDEC/NET0122_XXDec/XI39/XI23/MM0_d
+ N_XXDEC/XI39/NET22_XXDec/XI39/XI23/MM0_g
+ N_XXDEC/XI39/XI23/NET32_XXDec/XI39/XI23/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI24/MM0 N_XXDEC/NET190_XXDec/XI39/XI24/MM0_d
+ N_X_SEL_FF<3>_XXDec/XI39/XI24/MM0_g
+ N_XXDEC/XI39/XI24/NET32_XXDec/XI39/XI24/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI27/MM0 N_XXDEC/NET0130_XXDec/XI39/XI27/MM0_d
+ N_XXDEC/XI39/NET22_XXDec/XI39/XI27/MM0_g
+ N_XXDEC/XI39/XI27/NET32_XXDec/XI39/XI27/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI7/MM1 N_WL<63>_XXDec/XI36/XI7/MM1_d
+ N_XXDEC/NET0137_XXDec/XI36/XI7/MM1_g N_VSS_XXDec/XI36/XI7/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI7/MM1 N_WL<55>_XXDec/XI35/XI7/MM1_d
+ N_XXDEC/NET0137_XXDec/XI35/XI7/MM1_g N_VSS_XXDec/XI35/XI7/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI7/MM1 N_WL<47>_XXDec/XI34/XI7/MM1_d
+ N_XXDEC/NET0137_XXDec/XI34/XI7/MM1_g N_VSS_XXDec/XI34/XI7/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI7/MM1 N_WL<39>_XXDec/XI33/XI7/MM1_d
+ N_XXDEC/NET0137_XXDec/XI33/XI7/MM1_g N_VSS_XXDec/XI33/XI7/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI7/MM1 N_WL<31>_XXDec/XI32/XI7/MM1_d
+ N_XXDEC/NET0137_XXDec/XI32/XI7/MM1_g N_VSS_XXDec/XI32/XI7/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI7/MM1 N_WL<23>_XXDec/XI31/XI7/MM1_d
+ N_XXDEC/NET0137_XXDec/XI31/XI7/MM1_g N_VSS_XXDec/XI31/XI7/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI7/MM1 N_WL<15>_XXDec/XI30/XI7/MM1_d
+ N_XXDEC/NET0137_XXDec/XI30/XI7/MM1_g N_VSS_XXDec/XI30/XI7/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI7/MM1 N_WL<7>_XXDec/XI27/XI7/MM1_d
+ N_XXDEC/NET0137_XXDec/XI27/XI7/MM1_g N_VSS_XXDec/XI27/XI7/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI7/MM0 N_WL<63>_XXDec/XI36/XI7/MM0_d
+ N_XXDEC/NET0123_XXDec/XI36/XI7/MM0_g N_VSS_XXDec/XI36/XI7/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI7/MM0 N_WL<55>_XXDec/XI35/XI7/MM0_d
+ N_XXDEC/NET187_XXDec/XI35/XI7/MM0_g N_VSS_XXDec/XI35/XI7/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI7/MM0 N_WL<47>_XXDec/XI34/XI7/MM0_d
+ N_XXDEC/NET188_XXDec/XI34/XI7/MM0_g N_VSS_XXDec/XI34/XI7/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI7/MM0 N_WL<39>_XXDec/XI33/XI7/MM0_d
+ N_XXDEC/NET0122_XXDec/XI33/XI7/MM0_g N_VSS_XXDec/XI33/XI7/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI7/MM0 N_WL<31>_XXDec/XI32/XI7/MM0_d
+ N_XXDEC/NET190_XXDec/XI32/XI7/MM0_g N_VSS_XXDec/XI32/XI7/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI7/MM0 N_WL<23>_XXDec/XI31/XI7/MM0_d
+ N_XXDEC/NET0220_XXDec/XI31/XI7/MM0_g N_VSS_XXDec/XI31/XI7/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI7/MM0 N_WL<15>_XXDec/XI30/XI7/MM0_d
+ N_XXDEC/NET192_XXDec/XI30/XI7/MM0_g N_VSS_XXDec/XI30/XI7/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI7/MM0 N_WL<7>_XXDec/XI27/XI7/MM0_d
+ N_XXDEC/NET0130_XXDec/XI27/XI7/MM0_g N_VSS_XXDec/XI27/XI7/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI6/MM1 N_WL<62>_XXDec/XI36/XI6/MM1_d
+ N_XXDEC/NET0138_XXDec/XI36/XI6/MM1_g N_VSS_XXDec/XI36/XI6/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI6/MM1 N_WL<54>_XXDec/XI35/XI6/MM1_d
+ N_XXDEC/NET0138_XXDec/XI35/XI6/MM1_g N_VSS_XXDec/XI35/XI6/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI6/MM1 N_WL<46>_XXDec/XI34/XI6/MM1_d
+ N_XXDEC/NET0138_XXDec/XI34/XI6/MM1_g N_VSS_XXDec/XI34/XI6/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI6/MM1 N_WL<38>_XXDec/XI33/XI6/MM1_d
+ N_XXDEC/NET0138_XXDec/XI33/XI6/MM1_g N_VSS_XXDec/XI33/XI6/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI6/MM1 N_WL<30>_XXDec/XI32/XI6/MM1_d
+ N_XXDEC/NET0138_XXDec/XI32/XI6/MM1_g N_VSS_XXDec/XI32/XI6/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI6/MM1 N_WL<22>_XXDec/XI31/XI6/MM1_d
+ N_XXDEC/NET0138_XXDec/XI31/XI6/MM1_g N_VSS_XXDec/XI31/XI6/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI6/MM1 N_WL<14>_XXDec/XI30/XI6/MM1_d
+ N_XXDEC/NET0138_XXDec/XI30/XI6/MM1_g N_VSS_XXDec/XI30/XI6/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI6/MM1 N_WL<6>_XXDec/XI27/XI6/MM1_d
+ N_XXDEC/NET0138_XXDec/XI27/XI6/MM1_g N_VSS_XXDec/XI27/XI6/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI6/MM0 N_WL<62>_XXDec/XI36/XI6/MM0_d
+ N_XXDEC/NET0123_XXDec/XI36/XI6/MM0_g N_VSS_XXDec/XI36/XI6/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI6/MM0 N_WL<54>_XXDec/XI35/XI6/MM0_d
+ N_XXDEC/NET187_XXDec/XI35/XI6/MM0_g N_VSS_XXDec/XI35/XI6/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI6/MM0 N_WL<46>_XXDec/XI34/XI6/MM0_d
+ N_XXDEC/NET188_XXDec/XI34/XI6/MM0_g N_VSS_XXDec/XI34/XI6/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI6/MM0 N_WL<38>_XXDec/XI33/XI6/MM0_d
+ N_XXDEC/NET0122_XXDec/XI33/XI6/MM0_g N_VSS_XXDec/XI33/XI6/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI6/MM0 N_WL<30>_XXDec/XI32/XI6/MM0_d
+ N_XXDEC/NET190_XXDec/XI32/XI6/MM0_g N_VSS_XXDec/XI32/XI6/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI6/MM0 N_WL<22>_XXDec/XI31/XI6/MM0_d
+ N_XXDEC/NET0220_XXDec/XI31/XI6/MM0_g N_VSS_XXDec/XI31/XI6/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI6/MM0 N_WL<14>_XXDec/XI30/XI6/MM0_d
+ N_XXDEC/NET192_XXDec/XI30/XI6/MM0_g N_VSS_XXDec/XI30/XI6/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI6/MM0 N_WL<6>_XXDec/XI27/XI6/MM0_d
+ N_XXDEC/NET0130_XXDec/XI27/XI6/MM0_g N_VSS_XXDec/XI27/XI6/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI5/MM1 N_WL<61>_XXDec/XI36/XI5/MM1_d
+ N_XXDEC/NET0139_XXDec/XI36/XI5/MM1_g N_VSS_XXDec/XI36/XI5/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI5/MM1 N_WL<53>_XXDec/XI35/XI5/MM1_d
+ N_XXDEC/NET0139_XXDec/XI35/XI5/MM1_g N_VSS_XXDec/XI35/XI5/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI5/MM1 N_WL<45>_XXDec/XI34/XI5/MM1_d
+ N_XXDEC/NET0139_XXDec/XI34/XI5/MM1_g N_VSS_XXDec/XI34/XI5/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI5/MM1 N_WL<37>_XXDec/XI33/XI5/MM1_d
+ N_XXDEC/NET0139_XXDec/XI33/XI5/MM1_g N_VSS_XXDec/XI33/XI5/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI5/MM1 N_WL<29>_XXDec/XI32/XI5/MM1_d
+ N_XXDEC/NET0139_XXDec/XI32/XI5/MM1_g N_VSS_XXDec/XI32/XI5/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI5/MM1 N_WL<21>_XXDec/XI31/XI5/MM1_d
+ N_XXDEC/NET0139_XXDec/XI31/XI5/MM1_g N_VSS_XXDec/XI31/XI5/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI5/MM1 N_WL<13>_XXDec/XI30/XI5/MM1_d
+ N_XXDEC/NET0139_XXDec/XI30/XI5/MM1_g N_VSS_XXDec/XI30/XI5/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI5/MM1 N_WL<5>_XXDec/XI27/XI5/MM1_d
+ N_XXDEC/NET0139_XXDec/XI27/XI5/MM1_g N_VSS_XXDec/XI27/XI5/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI5/MM0 N_WL<61>_XXDec/XI36/XI5/MM0_d
+ N_XXDEC/NET0123_XXDec/XI36/XI5/MM0_g N_VSS_XXDec/XI36/XI5/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI5/MM0 N_WL<53>_XXDec/XI35/XI5/MM0_d
+ N_XXDEC/NET187_XXDec/XI35/XI5/MM0_g N_VSS_XXDec/XI35/XI5/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI5/MM0 N_WL<45>_XXDec/XI34/XI5/MM0_d
+ N_XXDEC/NET188_XXDec/XI34/XI5/MM0_g N_VSS_XXDec/XI34/XI5/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI5/MM0 N_WL<37>_XXDec/XI33/XI5/MM0_d
+ N_XXDEC/NET0122_XXDec/XI33/XI5/MM0_g N_VSS_XXDec/XI33/XI5/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI5/MM0 N_WL<29>_XXDec/XI32/XI5/MM0_d
+ N_XXDEC/NET190_XXDec/XI32/XI5/MM0_g N_VSS_XXDec/XI32/XI5/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI5/MM0 N_WL<21>_XXDec/XI31/XI5/MM0_d
+ N_XXDEC/NET0220_XXDec/XI31/XI5/MM0_g N_VSS_XXDec/XI31/XI5/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI5/MM0 N_WL<13>_XXDec/XI30/XI5/MM0_d
+ N_XXDEC/NET192_XXDec/XI30/XI5/MM0_g N_VSS_XXDec/XI30/XI5/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI5/MM0 N_WL<5>_XXDec/XI27/XI5/MM0_d
+ N_XXDEC/NET0130_XXDec/XI27/XI5/MM0_g N_VSS_XXDec/XI27/XI5/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI4/MM1 N_WL<60>_XXDec/XI36/XI4/MM1_d
+ N_XXDEC/NET0140_XXDec/XI36/XI4/MM1_g N_VSS_XXDec/XI36/XI4/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI4/MM1 N_WL<52>_XXDec/XI35/XI4/MM1_d
+ N_XXDEC/NET0140_XXDec/XI35/XI4/MM1_g N_VSS_XXDec/XI35/XI4/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI4/MM1 N_WL<44>_XXDec/XI34/XI4/MM1_d
+ N_XXDEC/NET0140_XXDec/XI34/XI4/MM1_g N_VSS_XXDec/XI34/XI4/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI4/MM1 N_WL<36>_XXDec/XI33/XI4/MM1_d
+ N_XXDEC/NET0140_XXDec/XI33/XI4/MM1_g N_VSS_XXDec/XI33/XI4/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI4/MM1 N_WL<28>_XXDec/XI32/XI4/MM1_d
+ N_XXDEC/NET0140_XXDec/XI32/XI4/MM1_g N_VSS_XXDec/XI32/XI4/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI4/MM1 N_WL<20>_XXDec/XI31/XI4/MM1_d
+ N_XXDEC/NET0140_XXDec/XI31/XI4/MM1_g N_VSS_XXDec/XI31/XI4/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI4/MM1 N_WL<12>_XXDec/XI30/XI4/MM1_d
+ N_XXDEC/NET0140_XXDec/XI30/XI4/MM1_g N_VSS_XXDec/XI30/XI4/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI4/MM1 N_WL<4>_XXDec/XI27/XI4/MM1_d
+ N_XXDEC/NET0140_XXDec/XI27/XI4/MM1_g N_VSS_XXDec/XI27/XI4/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI4/MM0 N_WL<60>_XXDec/XI36/XI4/MM0_d
+ N_XXDEC/NET0123_XXDec/XI36/XI4/MM0_g N_VSS_XXDec/XI36/XI4/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI4/MM0 N_WL<52>_XXDec/XI35/XI4/MM0_d
+ N_XXDEC/NET187_XXDec/XI35/XI4/MM0_g N_VSS_XXDec/XI35/XI4/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI4/MM0 N_WL<44>_XXDec/XI34/XI4/MM0_d
+ N_XXDEC/NET188_XXDec/XI34/XI4/MM0_g N_VSS_XXDec/XI34/XI4/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI4/MM0 N_WL<36>_XXDec/XI33/XI4/MM0_d
+ N_XXDEC/NET0122_XXDec/XI33/XI4/MM0_g N_VSS_XXDec/XI33/XI4/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI4/MM0 N_WL<28>_XXDec/XI32/XI4/MM0_d
+ N_XXDEC/NET190_XXDec/XI32/XI4/MM0_g N_VSS_XXDec/XI32/XI4/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI4/MM0 N_WL<20>_XXDec/XI31/XI4/MM0_d
+ N_XXDEC/NET0220_XXDec/XI31/XI4/MM0_g N_VSS_XXDec/XI31/XI4/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI4/MM0 N_WL<12>_XXDec/XI30/XI4/MM0_d
+ N_XXDEC/NET192_XXDec/XI30/XI4/MM0_g N_VSS_XXDec/XI30/XI4/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI4/MM0 N_WL<4>_XXDec/XI27/XI4/MM0_d
+ N_XXDEC/NET0130_XXDec/XI27/XI4/MM0_g N_VSS_XXDec/XI27/XI4/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI3/MM1 N_WL<59>_XXDec/XI36/XI3/MM1_d
+ N_XXDEC/NET0141_XXDec/XI36/XI3/MM1_g N_VSS_XXDec/XI36/XI3/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI3/MM1 N_WL<51>_XXDec/XI35/XI3/MM1_d
+ N_XXDEC/NET0141_XXDec/XI35/XI3/MM1_g N_VSS_XXDec/XI35/XI3/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI3/MM1 N_WL<43>_XXDec/XI34/XI3/MM1_d
+ N_XXDEC/NET0141_XXDec/XI34/XI3/MM1_g N_VSS_XXDec/XI34/XI3/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI3/MM1 N_WL<35>_XXDec/XI33/XI3/MM1_d
+ N_XXDEC/NET0141_XXDec/XI33/XI3/MM1_g N_VSS_XXDec/XI33/XI3/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI3/MM1 N_WL<27>_XXDec/XI32/XI3/MM1_d
+ N_XXDEC/NET0141_XXDec/XI32/XI3/MM1_g N_VSS_XXDec/XI32/XI3/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI3/MM1 N_WL<19>_XXDec/XI31/XI3/MM1_d
+ N_XXDEC/NET0141_XXDec/XI31/XI3/MM1_g N_VSS_XXDec/XI31/XI3/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI3/MM1 N_WL<11>_XXDec/XI30/XI3/MM1_d
+ N_XXDEC/NET0141_XXDec/XI30/XI3/MM1_g N_VSS_XXDec/XI30/XI3/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI3/MM1 N_WL<3>_XXDec/XI27/XI3/MM1_d
+ N_XXDEC/NET0141_XXDec/XI27/XI3/MM1_g N_VSS_XXDec/XI27/XI3/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI3/MM0 N_WL<59>_XXDec/XI36/XI3/MM0_d
+ N_XXDEC/NET0123_XXDec/XI36/XI3/MM0_g N_VSS_XXDec/XI36/XI3/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI3/MM0 N_WL<51>_XXDec/XI35/XI3/MM0_d
+ N_XXDEC/NET187_XXDec/XI35/XI3/MM0_g N_VSS_XXDec/XI35/XI3/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI3/MM0 N_WL<43>_XXDec/XI34/XI3/MM0_d
+ N_XXDEC/NET188_XXDec/XI34/XI3/MM0_g N_VSS_XXDec/XI34/XI3/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI3/MM0 N_WL<35>_XXDec/XI33/XI3/MM0_d
+ N_XXDEC/NET0122_XXDec/XI33/XI3/MM0_g N_VSS_XXDec/XI33/XI3/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI3/MM0 N_WL<27>_XXDec/XI32/XI3/MM0_d
+ N_XXDEC/NET190_XXDec/XI32/XI3/MM0_g N_VSS_XXDec/XI32/XI3/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI3/MM0 N_WL<19>_XXDec/XI31/XI3/MM0_d
+ N_XXDEC/NET0220_XXDec/XI31/XI3/MM0_g N_VSS_XXDec/XI31/XI3/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI3/MM0 N_WL<11>_XXDec/XI30/XI3/MM0_d
+ N_XXDEC/NET192_XXDec/XI30/XI3/MM0_g N_VSS_XXDec/XI30/XI3/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI3/MM0 N_WL<3>_XXDec/XI27/XI3/MM0_d
+ N_XXDEC/NET0130_XXDec/XI27/XI3/MM0_g N_VSS_XXDec/XI27/XI3/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI2/MM1 N_WL<58>_XXDec/XI36/XI2/MM1_d
+ N_XXDEC/NET0142_XXDec/XI36/XI2/MM1_g N_VSS_XXDec/XI36/XI2/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI2/MM1 N_WL<50>_XXDec/XI35/XI2/MM1_d
+ N_XXDEC/NET0142_XXDec/XI35/XI2/MM1_g N_VSS_XXDec/XI35/XI2/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI2/MM1 N_WL<42>_XXDec/XI34/XI2/MM1_d
+ N_XXDEC/NET0142_XXDec/XI34/XI2/MM1_g N_VSS_XXDec/XI34/XI2/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI2/MM1 N_WL<34>_XXDec/XI33/XI2/MM1_d
+ N_XXDEC/NET0142_XXDec/XI33/XI2/MM1_g N_VSS_XXDec/XI33/XI2/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI2/MM1 N_WL<26>_XXDec/XI32/XI2/MM1_d
+ N_XXDEC/NET0142_XXDec/XI32/XI2/MM1_g N_VSS_XXDec/XI32/XI2/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI2/MM1 N_WL<18>_XXDec/XI31/XI2/MM1_d
+ N_XXDEC/NET0142_XXDec/XI31/XI2/MM1_g N_VSS_XXDec/XI31/XI2/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI2/MM1 N_WL<10>_XXDec/XI30/XI2/MM1_d
+ N_XXDEC/NET0142_XXDec/XI30/XI2/MM1_g N_VSS_XXDec/XI30/XI2/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI2/MM1 N_WL<2>_XXDec/XI27/XI2/MM1_d
+ N_XXDEC/NET0142_XXDec/XI27/XI2/MM1_g N_VSS_XXDec/XI27/XI2/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI2/MM0 N_WL<58>_XXDec/XI36/XI2/MM0_d
+ N_XXDEC/NET0123_XXDec/XI36/XI2/MM0_g N_VSS_XXDec/XI36/XI2/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI2/MM0 N_WL<50>_XXDec/XI35/XI2/MM0_d
+ N_XXDEC/NET187_XXDec/XI35/XI2/MM0_g N_VSS_XXDec/XI35/XI2/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI2/MM0 N_WL<42>_XXDec/XI34/XI2/MM0_d
+ N_XXDEC/NET188_XXDec/XI34/XI2/MM0_g N_VSS_XXDec/XI34/XI2/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI2/MM0 N_WL<34>_XXDec/XI33/XI2/MM0_d
+ N_XXDEC/NET0122_XXDec/XI33/XI2/MM0_g N_VSS_XXDec/XI33/XI2/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI2/MM0 N_WL<26>_XXDec/XI32/XI2/MM0_d
+ N_XXDEC/NET190_XXDec/XI32/XI2/MM0_g N_VSS_XXDec/XI32/XI2/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI2/MM0 N_WL<18>_XXDec/XI31/XI2/MM0_d
+ N_XXDEC/NET0220_XXDec/XI31/XI2/MM0_g N_VSS_XXDec/XI31/XI2/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI2/MM0 N_WL<10>_XXDec/XI30/XI2/MM0_d
+ N_XXDEC/NET192_XXDec/XI30/XI2/MM0_g N_VSS_XXDec/XI30/XI2/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI2/MM0 N_WL<2>_XXDec/XI27/XI2/MM0_d
+ N_XXDEC/NET0130_XXDec/XI27/XI2/MM0_g N_VSS_XXDec/XI27/XI2/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI1/MM1 N_WL<57>_XXDec/XI36/XI1/MM1_d
+ N_XXDEC/NET0143_XXDec/XI36/XI1/MM1_g N_VSS_XXDec/XI36/XI1/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI1/MM1 N_WL<49>_XXDec/XI35/XI1/MM1_d
+ N_XXDEC/NET0143_XXDec/XI35/XI1/MM1_g N_VSS_XXDec/XI35/XI1/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI1/MM1 N_WL<41>_XXDec/XI34/XI1/MM1_d
+ N_XXDEC/NET0143_XXDec/XI34/XI1/MM1_g N_VSS_XXDec/XI34/XI1/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI1/MM1 N_WL<33>_XXDec/XI33/XI1/MM1_d
+ N_XXDEC/NET0143_XXDec/XI33/XI1/MM1_g N_VSS_XXDec/XI33/XI1/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI1/MM1 N_WL<25>_XXDec/XI32/XI1/MM1_d
+ N_XXDEC/NET0143_XXDec/XI32/XI1/MM1_g N_VSS_XXDec/XI32/XI1/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI1/MM1 N_WL<17>_XXDec/XI31/XI1/MM1_d
+ N_XXDEC/NET0143_XXDec/XI31/XI1/MM1_g N_VSS_XXDec/XI31/XI1/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI1/MM1 N_WL<9>_XXDec/XI30/XI1/MM1_d
+ N_XXDEC/NET0143_XXDec/XI30/XI1/MM1_g N_VSS_XXDec/XI30/XI1/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI1/MM1 N_WL<1>_XXDec/XI27/XI1/MM1_d
+ N_XXDEC/NET0143_XXDec/XI27/XI1/MM1_g N_VSS_XXDec/XI27/XI1/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI1/MM0 N_WL<57>_XXDec/XI36/XI1/MM0_d
+ N_XXDEC/NET0123_XXDec/XI36/XI1/MM0_g N_VSS_XXDec/XI36/XI1/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI1/MM0 N_WL<49>_XXDec/XI35/XI1/MM0_d
+ N_XXDEC/NET187_XXDec/XI35/XI1/MM0_g N_VSS_XXDec/XI35/XI1/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI1/MM0 N_WL<41>_XXDec/XI34/XI1/MM0_d
+ N_XXDEC/NET188_XXDec/XI34/XI1/MM0_g N_VSS_XXDec/XI34/XI1/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI1/MM0 N_WL<33>_XXDec/XI33/XI1/MM0_d
+ N_XXDEC/NET0122_XXDec/XI33/XI1/MM0_g N_VSS_XXDec/XI33/XI1/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI1/MM0 N_WL<25>_XXDec/XI32/XI1/MM0_d
+ N_XXDEC/NET190_XXDec/XI32/XI1/MM0_g N_VSS_XXDec/XI32/XI1/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI1/MM0 N_WL<17>_XXDec/XI31/XI1/MM0_d
+ N_XXDEC/NET0220_XXDec/XI31/XI1/MM0_g N_VSS_XXDec/XI31/XI1/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI1/MM0 N_WL<9>_XXDec/XI30/XI1/MM0_d
+ N_XXDEC/NET192_XXDec/XI30/XI1/MM0_g N_VSS_XXDec/XI30/XI1/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI1/MM0 N_WL<1>_XXDec/XI27/XI1/MM0_d
+ N_XXDEC/NET0130_XXDec/XI27/XI1/MM0_g N_VSS_XXDec/XI27/XI1/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI0/MM1 N_WL<56>_XXDec/XI36/XI0/MM1_d
+ N_XXDEC/NET0144_XXDec/XI36/XI0/MM1_g N_VSS_XXDec/XI36/XI0/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI0/MM1 N_WL<48>_XXDec/XI35/XI0/MM1_d
+ N_XXDEC/NET0144_XXDec/XI35/XI0/MM1_g N_VSS_XXDec/XI35/XI0/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI0/MM1 N_WL<40>_XXDec/XI34/XI0/MM1_d
+ N_XXDEC/NET0144_XXDec/XI34/XI0/MM1_g N_VSS_XXDec/XI34/XI0/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI0/MM1 N_WL<32>_XXDec/XI33/XI0/MM1_d
+ N_XXDEC/NET0144_XXDec/XI33/XI0/MM1_g N_VSS_XXDec/XI33/XI0/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI0/MM1 N_WL<24>_XXDec/XI32/XI0/MM1_d
+ N_XXDEC/NET0144_XXDec/XI32/XI0/MM1_g N_VSS_XXDec/XI32/XI0/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI0/MM1 N_WL<16>_XXDec/XI31/XI0/MM1_d
+ N_XXDEC/NET0144_XXDec/XI31/XI0/MM1_g N_VSS_XXDec/XI31/XI0/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI0/MM1 N_WL<8>_XXDec/XI30/XI0/MM1_d
+ N_XXDEC/NET0144_XXDec/XI30/XI0/MM1_g N_VSS_XXDec/XI30/XI0/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI0/MM1 N_WL<0>_XXDec/XI27/XI0/MM1_d
+ N_XXDEC/NET0144_XXDec/XI27/XI0/MM1_g N_VSS_XXDec/XI27/XI0/MM1_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI0/MM0 N_WL<56>_XXDec/XI36/XI0/MM0_d
+ N_XXDEC/NET0123_XXDec/XI36/XI0/MM0_g N_VSS_XXDec/XI36/XI0/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI0/MM0 N_WL<48>_XXDec/XI35/XI0/MM0_d
+ N_XXDEC/NET187_XXDec/XI35/XI0/MM0_g N_VSS_XXDec/XI35/XI0/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI0/MM0 N_WL<40>_XXDec/XI34/XI0/MM0_d
+ N_XXDEC/NET188_XXDec/XI34/XI0/MM0_g N_VSS_XXDec/XI34/XI0/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI0/MM0 N_WL<32>_XXDec/XI33/XI0/MM0_d
+ N_XXDEC/NET0122_XXDec/XI33/XI0/MM0_g N_VSS_XXDec/XI33/XI0/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI0/MM0 N_WL<24>_XXDec/XI32/XI0/MM0_d
+ N_XXDEC/NET190_XXDec/XI32/XI0/MM0_g N_VSS_XXDec/XI32/XI0/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI0/MM0 N_WL<16>_XXDec/XI31/XI0/MM0_d
+ N_XXDEC/NET0220_XXDec/XI31/XI0/MM0_g N_VSS_XXDec/XI31/XI0/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI0/MM0 N_WL<8>_XXDec/XI30/XI0/MM0_d
+ N_XXDEC/NET192_XXDec/XI30/XI0/MM0_g N_VSS_XXDec/XI30/XI0/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI0/MM0 N_WL<0>_XXDec/XI27/XI0/MM0_d
+ N_XXDEC/NET0130_XXDec/XI27/XI0/MM0_g N_VSS_XXDec/XI27/XI0/MM0_s
+ N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI17/MP N_XXDEC/XI40/NET22_XXDec/XI40/XI17/MP_d
+ N_X_SEL_FF<0>_XXDec/XI40/XI17/MP_g N_VDD_XXDec/XI40/XI17/MP_s
+ N_VDD_XXDec/XI40/XI17/MP_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXXDec/XI39/XI17/MP N_XXDEC/XI39/NET22_XXDec/XI39/XI17/MP_d
+ N_X_SEL_FF<3>_XXDec/XI39/XI17/MP_g N_VDD_XXDec/XI39/XI17/MP_s
+ N_VDD_XXDec/XI39/XI17/MP_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXXDec/XI40/XI18/MP N_XXDEC/XI40/NET18_XXDec/XI40/XI18/MP_d
+ N_X_SEL_FF<1>_XXDec/XI40/XI18/MP_g N_VDD_XXDec/XI40/XI18/MP_s
+ N_VDD_XXDec/XI40/XI18/MP_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXXDec/XI39/XI18/MP N_XXDEC/XI39/NET18_XXDec/XI39/XI18/MP_d
+ N_X_SEL_FF<4>_XXDec/XI39/XI18/MP_g N_VDD_XXDec/XI39/XI18/MP_s
+ N_VDD_XXDec/XI39/XI18/MP_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXXDec/XI40/XI19/MP N_XXDEC/XI40/NET14_XXDec/XI40/XI19/MP_d
+ N_X_SEL_FF<2>_XXDec/XI40/XI19/MP_g N_VDD_XXDec/XI40/XI19/MP_s
+ N_VDD_XXDec/XI40/XI19/MP_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXXDec/XI39/XI19/MP N_XXDEC/XI39/NET14_XXDec/XI39/XI19/MP_d
+ N_X_SEL_FF<5>_XXDec/XI39/XI19/MP_g N_VDD_XXDec/XI39/XI19/MP_s
+ N_VDD_XXDec/XI39/XI19/MP_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXXDec/XI40/XI26/MM7 N_XXDEC/NET0143_XXDec/XI40/XI26/MM7_d
+ N_WL_EN_XXDec/XI40/XI26/MM7_g N_VDD_XXDec/XI40/XI26/MM7_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI25/MM7 N_XXDEC/NET0142_XXDec/XI40/XI25/MM7_d
+ N_WL_EN_XXDec/XI40/XI25/MM7_g N_VDD_XXDec/XI40/XI25/MM7_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI22/MM7 N_XXDEC/NET0139_XXDec/XI40/XI22/MM7_d
+ N_WL_EN_XXDec/XI40/XI22/MM7_g N_VDD_XXDec/XI40/XI22/MM7_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI21/MM7 N_XXDEC/NET0138_XXDec/XI40/XI21/MM7_d
+ N_WL_EN_XXDec/XI40/XI21/MM7_g N_VDD_XXDec/XI40/XI21/MM7_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI21/MM7 N_XXDEC/NET187_XXDec/XI39/XI21/MM7_d
+ N_WL_EN_XXDec/XI39/XI21/MM7_g N_VDD_XXDec/XI39/XI21/MM7_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI22/MM7 N_XXDEC/NET188_XXDec/XI39/XI22/MM7_d
+ N_WL_EN_XXDec/XI39/XI22/MM7_g N_VDD_XXDec/XI39/XI22/MM7_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI25/MM7 N_XXDEC/NET0220_XXDec/XI39/XI25/MM7_d
+ N_WL_EN_XXDec/XI39/XI25/MM7_g N_VDD_XXDec/XI39/XI25/MM7_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI26/MM7 N_XXDEC/NET192_XXDec/XI39/XI26/MM7_d
+ N_WL_EN_XXDec/XI39/XI26/MM7_g N_VDD_XXDec/XI39/XI26/MM7_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI26/MM4 N_XXDEC/NET0143_XXDec/XI40/XI26/MM4_d
+ N_XXDEC/XI40/NET14_XXDec/XI40/XI26/MM4_g N_VDD_XXDec/XI40/XI26/MM4_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI25/MM4 N_XXDEC/NET0142_XXDec/XI40/XI25/MM4_d
+ N_XXDEC/XI40/NET14_XXDec/XI40/XI25/MM4_g N_VDD_XXDec/XI40/XI25/MM4_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI22/MM4 N_XXDEC/NET0139_XXDec/XI40/XI22/MM4_d
+ N_X_SEL_FF<2>_XXDec/XI40/XI22/MM4_g N_VDD_XXDec/XI40/XI22/MM4_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI21/MM4 N_XXDEC/NET0138_XXDec/XI40/XI21/MM4_d
+ N_X_SEL_FF<2>_XXDec/XI40/XI21/MM4_g N_VDD_XXDec/XI40/XI21/MM4_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI21/MM4 N_XXDEC/NET187_XXDec/XI39/XI21/MM4_d
+ N_X_SEL_FF<5>_XXDec/XI39/XI21/MM4_g N_VDD_XXDec/XI39/XI21/MM4_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI22/MM4 N_XXDEC/NET188_XXDec/XI39/XI22/MM4_d
+ N_X_SEL_FF<5>_XXDec/XI39/XI22/MM4_g N_VDD_XXDec/XI39/XI22/MM4_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI25/MM4 N_XXDEC/NET0220_XXDec/XI39/XI25/MM4_d
+ N_XXDEC/XI39/NET14_XXDec/XI39/XI25/MM4_g N_VDD_XXDec/XI39/XI25/MM4_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI26/MM4 N_XXDEC/NET192_XXDec/XI39/XI26/MM4_d
+ N_XXDEC/XI39/NET14_XXDec/XI39/XI26/MM4_g N_VDD_XXDec/XI39/XI26/MM4_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI26/MM5 N_XXDEC/NET0143_XXDec/XI40/XI26/MM5_d
+ N_XXDEC/XI40/NET18_XXDec/XI40/XI26/MM5_g N_VDD_XXDec/XI40/XI26/MM5_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI25/MM5 N_XXDEC/NET0142_XXDec/XI40/XI25/MM5_d
+ N_X_SEL_FF<1>_XXDec/XI40/XI25/MM5_g N_VDD_XXDec/XI40/XI25/MM5_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI22/MM5 N_XXDEC/NET0139_XXDec/XI40/XI22/MM5_d
+ N_XXDEC/XI40/NET18_XXDec/XI40/XI22/MM5_g N_VDD_XXDec/XI40/XI22/MM5_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI21/MM5 N_XXDEC/NET0138_XXDec/XI40/XI21/MM5_d
+ N_X_SEL_FF<1>_XXDec/XI40/XI21/MM5_g N_VDD_XXDec/XI40/XI21/MM5_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI21/MM5 N_XXDEC/NET187_XXDec/XI39/XI21/MM5_d
+ N_X_SEL_FF<4>_XXDec/XI39/XI21/MM5_g N_VDD_XXDec/XI39/XI21/MM5_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI22/MM5 N_XXDEC/NET188_XXDec/XI39/XI22/MM5_d
+ N_XXDEC/XI39/NET18_XXDec/XI39/XI22/MM5_g N_VDD_XXDec/XI39/XI22/MM5_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI25/MM5 N_XXDEC/NET0220_XXDec/XI39/XI25/MM5_d
+ N_X_SEL_FF<4>_XXDec/XI39/XI25/MM5_g N_VDD_XXDec/XI39/XI25/MM5_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI26/MM5 N_XXDEC/NET192_XXDec/XI39/XI26/MM5_d
+ N_XXDEC/XI39/NET18_XXDec/XI39/XI26/MM5_g N_VDD_XXDec/XI39/XI26/MM5_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI26/MM6 N_XXDEC/NET0143_XXDec/XI40/XI26/MM6_d
+ N_X_SEL_FF<0>_XXDec/XI40/XI26/MM6_g N_VDD_XXDec/XI40/XI26/MM6_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI25/MM6 N_XXDEC/NET0142_XXDec/XI40/XI25/MM6_d
+ N_XXDEC/XI40/NET22_XXDec/XI40/XI25/MM6_g N_VDD_XXDec/XI40/XI25/MM6_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI22/MM6 N_XXDEC/NET0139_XXDec/XI40/XI22/MM6_d
+ N_X_SEL_FF<0>_XXDec/XI40/XI22/MM6_g N_VDD_XXDec/XI40/XI22/MM6_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI21/MM6 N_XXDEC/NET0138_XXDec/XI40/XI21/MM6_d
+ N_XXDEC/XI40/NET22_XXDec/XI40/XI21/MM6_g N_VDD_XXDec/XI40/XI21/MM6_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI21/MM6 N_XXDEC/NET187_XXDec/XI39/XI21/MM6_d
+ N_XXDEC/XI39/NET22_XXDec/XI39/XI21/MM6_g N_VDD_XXDec/XI39/XI21/MM6_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI22/MM6 N_XXDEC/NET188_XXDec/XI39/XI22/MM6_d
+ N_X_SEL_FF<3>_XXDec/XI39/XI22/MM6_g N_VDD_XXDec/XI39/XI22/MM6_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI25/MM6 N_XXDEC/NET0220_XXDec/XI39/XI25/MM6_d
+ N_XXDEC/XI39/NET22_XXDec/XI39/XI25/MM6_g N_VDD_XXDec/XI39/XI25/MM6_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI26/MM6 N_XXDEC/NET192_XXDec/XI39/XI26/MM6_d
+ N_X_SEL_FF<3>_XXDec/XI39/XI26/MM6_g N_VDD_XXDec/XI39/XI26/MM6_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI27/MM7 N_XXDEC/NET0144_XXDec/XI40/XI27/MM7_d
+ N_WL_EN_XXDec/XI40/XI27/MM7_g N_VDD_XXDec/XI40/XI27/MM7_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI24/MM7 N_XXDEC/NET0141_XXDec/XI40/XI24/MM7_d
+ N_WL_EN_XXDec/XI40/XI24/MM7_g N_VDD_XXDec/XI40/XI24/MM7_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI23/MM7 N_XXDEC/NET0140_XXDec/XI40/XI23/MM7_d
+ N_WL_EN_XXDec/XI40/XI23/MM7_g N_VDD_XXDec/XI40/XI23/MM7_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI20/MM7 N_XXDEC/NET0137_XXDec/XI40/XI20/MM7_d
+ N_WL_EN_XXDec/XI40/XI20/MM7_g N_VDD_XXDec/XI40/XI20/MM7_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI20/MM7 N_XXDEC/NET0123_XXDec/XI39/XI20/MM7_d
+ N_WL_EN_XXDec/XI39/XI20/MM7_g N_VDD_XXDec/XI39/XI20/MM7_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI23/MM7 N_XXDEC/NET0122_XXDec/XI39/XI23/MM7_d
+ N_WL_EN_XXDec/XI39/XI23/MM7_g N_VDD_XXDec/XI39/XI23/MM7_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI24/MM7 N_XXDEC/NET190_XXDec/XI39/XI24/MM7_d
+ N_WL_EN_XXDec/XI39/XI24/MM7_g N_VDD_XXDec/XI39/XI24/MM7_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI27/MM7 N_XXDEC/NET0130_XXDec/XI39/XI27/MM7_d
+ N_WL_EN_XXDec/XI39/XI27/MM7_g N_VDD_XXDec/XI39/XI27/MM7_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI27/MM4 N_XXDEC/NET0144_XXDec/XI40/XI27/MM4_d
+ N_XXDEC/XI40/NET14_XXDec/XI40/XI27/MM4_g N_VDD_XXDec/XI40/XI27/MM4_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI24/MM4 N_XXDEC/NET0141_XXDec/XI40/XI24/MM4_d
+ N_XXDEC/XI40/NET14_XXDec/XI40/XI24/MM4_g N_VDD_XXDec/XI40/XI24/MM4_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI23/MM4 N_XXDEC/NET0140_XXDec/XI40/XI23/MM4_d
+ N_X_SEL_FF<2>_XXDec/XI40/XI23/MM4_g N_VDD_XXDec/XI40/XI23/MM4_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI20/MM4 N_XXDEC/NET0137_XXDec/XI40/XI20/MM4_d
+ N_X_SEL_FF<2>_XXDec/XI40/XI20/MM4_g N_VDD_XXDec/XI40/XI20/MM4_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI20/MM4 N_XXDEC/NET0123_XXDec/XI39/XI20/MM4_d
+ N_X_SEL_FF<5>_XXDec/XI39/XI20/MM4_g N_VDD_XXDec/XI39/XI20/MM4_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI23/MM4 N_XXDEC/NET0122_XXDec/XI39/XI23/MM4_d
+ N_X_SEL_FF<5>_XXDec/XI39/XI23/MM4_g N_VDD_XXDec/XI39/XI23/MM4_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI24/MM4 N_XXDEC/NET190_XXDec/XI39/XI24/MM4_d
+ N_XXDEC/XI39/NET14_XXDec/XI39/XI24/MM4_g N_VDD_XXDec/XI39/XI24/MM4_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI27/MM4 N_XXDEC/NET0130_XXDec/XI39/XI27/MM4_d
+ N_XXDEC/XI39/NET14_XXDec/XI39/XI27/MM4_g N_VDD_XXDec/XI39/XI27/MM4_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI27/MM5 N_XXDEC/NET0144_XXDec/XI40/XI27/MM5_d
+ N_XXDEC/XI40/NET18_XXDec/XI40/XI27/MM5_g N_VDD_XXDec/XI40/XI27/MM5_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI24/MM5 N_XXDEC/NET0141_XXDec/XI40/XI24/MM5_d
+ N_X_SEL_FF<1>_XXDec/XI40/XI24/MM5_g N_VDD_XXDec/XI40/XI24/MM5_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI23/MM5 N_XXDEC/NET0140_XXDec/XI40/XI23/MM5_d
+ N_XXDEC/XI40/NET18_XXDec/XI40/XI23/MM5_g N_VDD_XXDec/XI40/XI23/MM5_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI20/MM5 N_XXDEC/NET0137_XXDec/XI40/XI20/MM5_d
+ N_X_SEL_FF<1>_XXDec/XI40/XI20/MM5_g N_VDD_XXDec/XI40/XI20/MM5_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI20/MM5 N_XXDEC/NET0123_XXDec/XI39/XI20/MM5_d
+ N_X_SEL_FF<4>_XXDec/XI39/XI20/MM5_g N_VDD_XXDec/XI39/XI20/MM5_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI23/MM5 N_XXDEC/NET0122_XXDec/XI39/XI23/MM5_d
+ N_XXDEC/XI39/NET18_XXDec/XI39/XI23/MM5_g N_VDD_XXDec/XI39/XI23/MM5_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI24/MM5 N_XXDEC/NET190_XXDec/XI39/XI24/MM5_d
+ N_X_SEL_FF<4>_XXDec/XI39/XI24/MM5_g N_VDD_XXDec/XI39/XI24/MM5_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI39/XI27/MM5 N_XXDEC/NET0130_XXDec/XI39/XI27/MM5_d
+ N_XXDEC/XI39/NET18_XXDec/XI39/XI27/MM5_g N_VDD_XXDec/XI39/XI27/MM5_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13
+ PD=5.1e-07 PS=5.1e-07
mXXDec/XI40/XI27/MM6 N_XXDEC/NET0144_XXDec/XI40/XI27/MM6_d
+ N_XXDEC/XI40/NET22_XXDec/XI40/XI27/MM6_g N_VDD_XXDec/XI40/XI27/MM6_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI24/MM6 N_XXDEC/NET0141_XXDec/XI40/XI24/MM6_d
+ N_X_SEL_FF<0>_XXDec/XI40/XI24/MM6_g N_VDD_XXDec/XI40/XI24/MM6_s
+ N_VDD_XXDec/XI40/XI26/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI23/MM6 N_XXDEC/NET0140_XXDec/XI40/XI23/MM6_d
+ N_XXDEC/XI40/NET22_XXDec/XI40/XI23/MM6_g N_VDD_XXDec/XI40/XI23/MM6_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI40/XI20/MM6 N_XXDEC/NET0137_XXDec/XI40/XI20/MM6_d
+ N_X_SEL_FF<0>_XXDec/XI40/XI20/MM6_g N_VDD_XXDec/XI40/XI20/MM6_s
+ N_VDD_XXDec/XI40/XI22/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI20/MM6 N_XXDEC/NET0123_XXDec/XI39/XI20/MM6_d
+ N_X_SEL_FF<3>_XXDec/XI39/XI20/MM6_g N_VDD_XXDec/XI39/XI20/MM6_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI23/MM6 N_XXDEC/NET0122_XXDec/XI39/XI23/MM6_d
+ N_XXDEC/XI39/NET22_XXDec/XI39/XI23/MM6_g N_VDD_XXDec/XI39/XI23/MM6_s
+ N_VDD_XXDec/XI39/XI21/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI24/MM6 N_XXDEC/NET190_XXDec/XI39/XI24/MM6_d
+ N_X_SEL_FF<3>_XXDec/XI39/XI24/MM6_g N_VDD_XXDec/XI39/XI24/MM6_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI39/XI27/MM6 N_XXDEC/NET0130_XXDec/XI39/XI27/MM6_d
+ N_XXDEC/XI39/NET22_XXDec/XI39/XI27/MM6_g N_VDD_XXDec/XI39/XI27/MM6_s
+ N_VDD_XXDec/XI39/XI25/MM7_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13
+ PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI7/MM2 N_XXDEC/XI36/XI7/NET13_XXDec/XI36/XI7/MM2_d
+ N_XXDEC/NET0137_XXDec/XI36/XI7/MM2_g N_VDD_XXDec/XI36/XI7/MM2_s
+ N_VDD_XXDec/XI36/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI35/XI7/MM2 N_XXDEC/XI35/XI7/NET13_XXDec/XI35/XI7/MM2_d
+ N_XXDEC/NET0137_XXDec/XI35/XI7/MM2_g N_VDD_XXDec/XI35/XI7/MM2_s
+ N_VDD_XXDec/XI35/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI34/XI7/MM2 N_XXDEC/XI34/XI7/NET13_XXDec/XI34/XI7/MM2_d
+ N_XXDEC/NET0137_XXDec/XI34/XI7/MM2_g N_VDD_XXDec/XI34/XI7/MM2_s
+ N_VDD_XXDec/XI34/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI33/XI7/MM2 N_XXDEC/XI33/XI7/NET13_XXDec/XI33/XI7/MM2_d
+ N_XXDEC/NET0137_XXDec/XI33/XI7/MM2_g N_VDD_XXDec/XI33/XI7/MM2_s
+ N_VDD_XXDec/XI33/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI32/XI7/MM2 N_XXDEC/XI32/XI7/NET13_XXDec/XI32/XI7/MM2_d
+ N_XXDEC/NET0137_XXDec/XI32/XI7/MM2_g N_VDD_XXDec/XI32/XI7/MM2_s
+ N_VDD_XXDec/XI32/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI31/XI7/MM2 N_XXDEC/XI31/XI7/NET13_XXDec/XI31/XI7/MM2_d
+ N_XXDEC/NET0137_XXDec/XI31/XI7/MM2_g N_VDD_XXDec/XI31/XI7/MM2_s
+ N_VDD_XXDec/XI31/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI30/XI7/MM2 N_XXDEC/XI30/XI7/NET13_XXDec/XI30/XI7/MM2_d
+ N_XXDEC/NET0137_XXDec/XI30/XI7/MM2_g N_VDD_XXDec/XI30/XI7/MM2_s
+ N_VDD_XXDec/XI30/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI27/XI7/MM2 N_XXDEC/XI27/XI7/NET13_XXDec/XI27/XI7/MM2_d
+ N_XXDEC/NET0137_XXDec/XI27/XI7/MM2_g N_VDD_XXDec/XI27/XI7/MM2_s
+ N_VDD_XXDec/XI27/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI36/XI7/MM3 N_WL<63>_XXDec/XI36/XI7/MM3_d
+ N_XXDEC/NET0123_XXDec/XI36/XI7/MM3_g
+ N_XXDEC/XI36/XI7/NET13_XXDec/XI36/XI7/MM3_s N_VDD_XXDec/XI36/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI7/MM3 N_WL<55>_XXDec/XI35/XI7/MM3_d
+ N_XXDEC/NET187_XXDec/XI35/XI7/MM3_g
+ N_XXDEC/XI35/XI7/NET13_XXDec/XI35/XI7/MM3_s N_VDD_XXDec/XI35/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI7/MM3 N_WL<47>_XXDec/XI34/XI7/MM3_d
+ N_XXDEC/NET188_XXDec/XI34/XI7/MM3_g
+ N_XXDEC/XI34/XI7/NET13_XXDec/XI34/XI7/MM3_s N_VDD_XXDec/XI34/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI7/MM3 N_WL<39>_XXDec/XI33/XI7/MM3_d
+ N_XXDEC/NET0122_XXDec/XI33/XI7/MM3_g
+ N_XXDEC/XI33/XI7/NET13_XXDec/XI33/XI7/MM3_s N_VDD_XXDec/XI33/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI7/MM3 N_WL<31>_XXDec/XI32/XI7/MM3_d
+ N_XXDEC/NET190_XXDec/XI32/XI7/MM3_g
+ N_XXDEC/XI32/XI7/NET13_XXDec/XI32/XI7/MM3_s N_VDD_XXDec/XI32/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI7/MM3 N_WL<23>_XXDec/XI31/XI7/MM3_d
+ N_XXDEC/NET0220_XXDec/XI31/XI7/MM3_g
+ N_XXDEC/XI31/XI7/NET13_XXDec/XI31/XI7/MM3_s N_VDD_XXDec/XI31/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI7/MM3 N_WL<15>_XXDec/XI30/XI7/MM3_d
+ N_XXDEC/NET192_XXDec/XI30/XI7/MM3_g
+ N_XXDEC/XI30/XI7/NET13_XXDec/XI30/XI7/MM3_s N_VDD_XXDec/XI30/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI7/MM3 N_WL<7>_XXDec/XI27/XI7/MM3_d
+ N_XXDEC/NET0130_XXDec/XI27/XI7/MM3_g
+ N_XXDEC/XI27/XI7/NET13_XXDec/XI27/XI7/MM3_s N_VDD_XXDec/XI27/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI6/MM2 N_XXDEC/XI36/XI6/NET13_XXDec/XI36/XI6/MM2_d
+ N_XXDEC/NET0138_XXDec/XI36/XI6/MM2_g N_VDD_XXDec/XI36/XI6/MM2_s
+ N_VDD_XXDec/XI36/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI35/XI6/MM2 N_XXDEC/XI35/XI6/NET13_XXDec/XI35/XI6/MM2_d
+ N_XXDEC/NET0138_XXDec/XI35/XI6/MM2_g N_VDD_XXDec/XI35/XI6/MM2_s
+ N_VDD_XXDec/XI35/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI34/XI6/MM2 N_XXDEC/XI34/XI6/NET13_XXDec/XI34/XI6/MM2_d
+ N_XXDEC/NET0138_XXDec/XI34/XI6/MM2_g N_VDD_XXDec/XI34/XI6/MM2_s
+ N_VDD_XXDec/XI34/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI33/XI6/MM2 N_XXDEC/XI33/XI6/NET13_XXDec/XI33/XI6/MM2_d
+ N_XXDEC/NET0138_XXDec/XI33/XI6/MM2_g N_VDD_XXDec/XI33/XI6/MM2_s
+ N_VDD_XXDec/XI33/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI32/XI6/MM2 N_XXDEC/XI32/XI6/NET13_XXDec/XI32/XI6/MM2_d
+ N_XXDEC/NET0138_XXDec/XI32/XI6/MM2_g N_VDD_XXDec/XI32/XI6/MM2_s
+ N_VDD_XXDec/XI32/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI31/XI6/MM2 N_XXDEC/XI31/XI6/NET13_XXDec/XI31/XI6/MM2_d
+ N_XXDEC/NET0138_XXDec/XI31/XI6/MM2_g N_VDD_XXDec/XI31/XI6/MM2_s
+ N_VDD_XXDec/XI31/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI30/XI6/MM2 N_XXDEC/XI30/XI6/NET13_XXDec/XI30/XI6/MM2_d
+ N_XXDEC/NET0138_XXDec/XI30/XI6/MM2_g N_VDD_XXDec/XI30/XI6/MM2_s
+ N_VDD_XXDec/XI30/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI27/XI6/MM2 N_XXDEC/XI27/XI6/NET13_XXDec/XI27/XI6/MM2_d
+ N_XXDEC/NET0138_XXDec/XI27/XI6/MM2_g N_VDD_XXDec/XI27/XI6/MM2_s
+ N_VDD_XXDec/XI27/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI36/XI6/MM3 N_WL<62>_XXDec/XI36/XI6/MM3_d
+ N_XXDEC/NET0123_XXDec/XI36/XI6/MM3_g
+ N_XXDEC/XI36/XI6/NET13_XXDec/XI36/XI6/MM3_s N_VDD_XXDec/XI36/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI6/MM3 N_WL<54>_XXDec/XI35/XI6/MM3_d
+ N_XXDEC/NET187_XXDec/XI35/XI6/MM3_g
+ N_XXDEC/XI35/XI6/NET13_XXDec/XI35/XI6/MM3_s N_VDD_XXDec/XI35/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI6/MM3 N_WL<46>_XXDec/XI34/XI6/MM3_d
+ N_XXDEC/NET188_XXDec/XI34/XI6/MM3_g
+ N_XXDEC/XI34/XI6/NET13_XXDec/XI34/XI6/MM3_s N_VDD_XXDec/XI34/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI6/MM3 N_WL<38>_XXDec/XI33/XI6/MM3_d
+ N_XXDEC/NET0122_XXDec/XI33/XI6/MM3_g
+ N_XXDEC/XI33/XI6/NET13_XXDec/XI33/XI6/MM3_s N_VDD_XXDec/XI33/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI6/MM3 N_WL<30>_XXDec/XI32/XI6/MM3_d
+ N_XXDEC/NET190_XXDec/XI32/XI6/MM3_g
+ N_XXDEC/XI32/XI6/NET13_XXDec/XI32/XI6/MM3_s N_VDD_XXDec/XI32/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI6/MM3 N_WL<22>_XXDec/XI31/XI6/MM3_d
+ N_XXDEC/NET0220_XXDec/XI31/XI6/MM3_g
+ N_XXDEC/XI31/XI6/NET13_XXDec/XI31/XI6/MM3_s N_VDD_XXDec/XI31/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI6/MM3 N_WL<14>_XXDec/XI30/XI6/MM3_d
+ N_XXDEC/NET192_XXDec/XI30/XI6/MM3_g
+ N_XXDEC/XI30/XI6/NET13_XXDec/XI30/XI6/MM3_s N_VDD_XXDec/XI30/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI6/MM3 N_WL<6>_XXDec/XI27/XI6/MM3_d
+ N_XXDEC/NET0130_XXDec/XI27/XI6/MM3_g
+ N_XXDEC/XI27/XI6/NET13_XXDec/XI27/XI6/MM3_s N_VDD_XXDec/XI27/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI5/MM2 N_XXDEC/XI36/XI5/NET13_XXDec/XI36/XI5/MM2_d
+ N_XXDEC/NET0139_XXDec/XI36/XI5/MM2_g N_VDD_XXDec/XI36/XI5/MM2_s
+ N_VDD_XXDec/XI36/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI35/XI5/MM2 N_XXDEC/XI35/XI5/NET13_XXDec/XI35/XI5/MM2_d
+ N_XXDEC/NET0139_XXDec/XI35/XI5/MM2_g N_VDD_XXDec/XI35/XI5/MM2_s
+ N_VDD_XXDec/XI35/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI34/XI5/MM2 N_XXDEC/XI34/XI5/NET13_XXDec/XI34/XI5/MM2_d
+ N_XXDEC/NET0139_XXDec/XI34/XI5/MM2_g N_VDD_XXDec/XI34/XI5/MM2_s
+ N_VDD_XXDec/XI34/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI33/XI5/MM2 N_XXDEC/XI33/XI5/NET13_XXDec/XI33/XI5/MM2_d
+ N_XXDEC/NET0139_XXDec/XI33/XI5/MM2_g N_VDD_XXDec/XI33/XI5/MM2_s
+ N_VDD_XXDec/XI33/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI32/XI5/MM2 N_XXDEC/XI32/XI5/NET13_XXDec/XI32/XI5/MM2_d
+ N_XXDEC/NET0139_XXDec/XI32/XI5/MM2_g N_VDD_XXDec/XI32/XI5/MM2_s
+ N_VDD_XXDec/XI32/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI31/XI5/MM2 N_XXDEC/XI31/XI5/NET13_XXDec/XI31/XI5/MM2_d
+ N_XXDEC/NET0139_XXDec/XI31/XI5/MM2_g N_VDD_XXDec/XI31/XI5/MM2_s
+ N_VDD_XXDec/XI31/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI30/XI5/MM2 N_XXDEC/XI30/XI5/NET13_XXDec/XI30/XI5/MM2_d
+ N_XXDEC/NET0139_XXDec/XI30/XI5/MM2_g N_VDD_XXDec/XI30/XI5/MM2_s
+ N_VDD_XXDec/XI30/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI27/XI5/MM2 N_XXDEC/XI27/XI5/NET13_XXDec/XI27/XI5/MM2_d
+ N_XXDEC/NET0139_XXDec/XI27/XI5/MM2_g N_VDD_XXDec/XI27/XI5/MM2_s
+ N_VDD_XXDec/XI27/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI36/XI5/MM3 N_WL<61>_XXDec/XI36/XI5/MM3_d
+ N_XXDEC/NET0123_XXDec/XI36/XI5/MM3_g
+ N_XXDEC/XI36/XI5/NET13_XXDec/XI36/XI5/MM3_s N_VDD_XXDec/XI36/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI5/MM3 N_WL<53>_XXDec/XI35/XI5/MM3_d
+ N_XXDEC/NET187_XXDec/XI35/XI5/MM3_g
+ N_XXDEC/XI35/XI5/NET13_XXDec/XI35/XI5/MM3_s N_VDD_XXDec/XI35/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI5/MM3 N_WL<45>_XXDec/XI34/XI5/MM3_d
+ N_XXDEC/NET188_XXDec/XI34/XI5/MM3_g
+ N_XXDEC/XI34/XI5/NET13_XXDec/XI34/XI5/MM3_s N_VDD_XXDec/XI34/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI5/MM3 N_WL<37>_XXDec/XI33/XI5/MM3_d
+ N_XXDEC/NET0122_XXDec/XI33/XI5/MM3_g
+ N_XXDEC/XI33/XI5/NET13_XXDec/XI33/XI5/MM3_s N_VDD_XXDec/XI33/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI5/MM3 N_WL<29>_XXDec/XI32/XI5/MM3_d
+ N_XXDEC/NET190_XXDec/XI32/XI5/MM3_g
+ N_XXDEC/XI32/XI5/NET13_XXDec/XI32/XI5/MM3_s N_VDD_XXDec/XI32/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI5/MM3 N_WL<21>_XXDec/XI31/XI5/MM3_d
+ N_XXDEC/NET0220_XXDec/XI31/XI5/MM3_g
+ N_XXDEC/XI31/XI5/NET13_XXDec/XI31/XI5/MM3_s N_VDD_XXDec/XI31/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI5/MM3 N_WL<13>_XXDec/XI30/XI5/MM3_d
+ N_XXDEC/NET192_XXDec/XI30/XI5/MM3_g
+ N_XXDEC/XI30/XI5/NET13_XXDec/XI30/XI5/MM3_s N_VDD_XXDec/XI30/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI5/MM3 N_WL<5>_XXDec/XI27/XI5/MM3_d
+ N_XXDEC/NET0130_XXDec/XI27/XI5/MM3_g
+ N_XXDEC/XI27/XI5/NET13_XXDec/XI27/XI5/MM3_s N_VDD_XXDec/XI27/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI4/MM2 N_XXDEC/XI36/XI4/NET13_XXDec/XI36/XI4/MM2_d
+ N_XXDEC/NET0140_XXDec/XI36/XI4/MM2_g N_VDD_XXDec/XI36/XI4/MM2_s
+ N_VDD_XXDec/XI36/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI35/XI4/MM2 N_XXDEC/XI35/XI4/NET13_XXDec/XI35/XI4/MM2_d
+ N_XXDEC/NET0140_XXDec/XI35/XI4/MM2_g N_VDD_XXDec/XI35/XI4/MM2_s
+ N_VDD_XXDec/XI35/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI34/XI4/MM2 N_XXDEC/XI34/XI4/NET13_XXDec/XI34/XI4/MM2_d
+ N_XXDEC/NET0140_XXDec/XI34/XI4/MM2_g N_VDD_XXDec/XI34/XI4/MM2_s
+ N_VDD_XXDec/XI34/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI33/XI4/MM2 N_XXDEC/XI33/XI4/NET13_XXDec/XI33/XI4/MM2_d
+ N_XXDEC/NET0140_XXDec/XI33/XI4/MM2_g N_VDD_XXDec/XI33/XI4/MM2_s
+ N_VDD_XXDec/XI33/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI32/XI4/MM2 N_XXDEC/XI32/XI4/NET13_XXDec/XI32/XI4/MM2_d
+ N_XXDEC/NET0140_XXDec/XI32/XI4/MM2_g N_VDD_XXDec/XI32/XI4/MM2_s
+ N_VDD_XXDec/XI32/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI31/XI4/MM2 N_XXDEC/XI31/XI4/NET13_XXDec/XI31/XI4/MM2_d
+ N_XXDEC/NET0140_XXDec/XI31/XI4/MM2_g N_VDD_XXDec/XI31/XI4/MM2_s
+ N_VDD_XXDec/XI31/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI30/XI4/MM2 N_XXDEC/XI30/XI4/NET13_XXDec/XI30/XI4/MM2_d
+ N_XXDEC/NET0140_XXDec/XI30/XI4/MM2_g N_VDD_XXDec/XI30/XI4/MM2_s
+ N_VDD_XXDec/XI30/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI27/XI4/MM2 N_XXDEC/XI27/XI4/NET13_XXDec/XI27/XI4/MM2_d
+ N_XXDEC/NET0140_XXDec/XI27/XI4/MM2_g N_VDD_XXDec/XI27/XI4/MM2_s
+ N_VDD_XXDec/XI27/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI36/XI4/MM3 N_WL<60>_XXDec/XI36/XI4/MM3_d
+ N_XXDEC/NET0123_XXDec/XI36/XI4/MM3_g
+ N_XXDEC/XI36/XI4/NET13_XXDec/XI36/XI4/MM3_s N_VDD_XXDec/XI36/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI4/MM3 N_WL<52>_XXDec/XI35/XI4/MM3_d
+ N_XXDEC/NET187_XXDec/XI35/XI4/MM3_g
+ N_XXDEC/XI35/XI4/NET13_XXDec/XI35/XI4/MM3_s N_VDD_XXDec/XI35/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI4/MM3 N_WL<44>_XXDec/XI34/XI4/MM3_d
+ N_XXDEC/NET188_XXDec/XI34/XI4/MM3_g
+ N_XXDEC/XI34/XI4/NET13_XXDec/XI34/XI4/MM3_s N_VDD_XXDec/XI34/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI4/MM3 N_WL<36>_XXDec/XI33/XI4/MM3_d
+ N_XXDEC/NET0122_XXDec/XI33/XI4/MM3_g
+ N_XXDEC/XI33/XI4/NET13_XXDec/XI33/XI4/MM3_s N_VDD_XXDec/XI33/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI4/MM3 N_WL<28>_XXDec/XI32/XI4/MM3_d
+ N_XXDEC/NET190_XXDec/XI32/XI4/MM3_g
+ N_XXDEC/XI32/XI4/NET13_XXDec/XI32/XI4/MM3_s N_VDD_XXDec/XI32/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI4/MM3 N_WL<20>_XXDec/XI31/XI4/MM3_d
+ N_XXDEC/NET0220_XXDec/XI31/XI4/MM3_g
+ N_XXDEC/XI31/XI4/NET13_XXDec/XI31/XI4/MM3_s N_VDD_XXDec/XI31/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI4/MM3 N_WL<12>_XXDec/XI30/XI4/MM3_d
+ N_XXDEC/NET192_XXDec/XI30/XI4/MM3_g
+ N_XXDEC/XI30/XI4/NET13_XXDec/XI30/XI4/MM3_s N_VDD_XXDec/XI30/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI4/MM3 N_WL<4>_XXDec/XI27/XI4/MM3_d
+ N_XXDEC/NET0130_XXDec/XI27/XI4/MM3_g
+ N_XXDEC/XI27/XI4/NET13_XXDec/XI27/XI4/MM3_s N_VDD_XXDec/XI27/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI3/MM2 N_XXDEC/XI36/XI3/NET13_XXDec/XI36/XI3/MM2_d
+ N_XXDEC/NET0141_XXDec/XI36/XI3/MM2_g N_VDD_XXDec/XI36/XI3/MM2_s
+ N_VDD_XXDec/XI36/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI35/XI3/MM2 N_XXDEC/XI35/XI3/NET13_XXDec/XI35/XI3/MM2_d
+ N_XXDEC/NET0141_XXDec/XI35/XI3/MM2_g N_VDD_XXDec/XI35/XI3/MM2_s
+ N_VDD_XXDec/XI35/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI34/XI3/MM2 N_XXDEC/XI34/XI3/NET13_XXDec/XI34/XI3/MM2_d
+ N_XXDEC/NET0141_XXDec/XI34/XI3/MM2_g N_VDD_XXDec/XI34/XI3/MM2_s
+ N_VDD_XXDec/XI34/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI33/XI3/MM2 N_XXDEC/XI33/XI3/NET13_XXDec/XI33/XI3/MM2_d
+ N_XXDEC/NET0141_XXDec/XI33/XI3/MM2_g N_VDD_XXDec/XI33/XI3/MM2_s
+ N_VDD_XXDec/XI33/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI32/XI3/MM2 N_XXDEC/XI32/XI3/NET13_XXDec/XI32/XI3/MM2_d
+ N_XXDEC/NET0141_XXDec/XI32/XI3/MM2_g N_VDD_XXDec/XI32/XI3/MM2_s
+ N_VDD_XXDec/XI32/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI31/XI3/MM2 N_XXDEC/XI31/XI3/NET13_XXDec/XI31/XI3/MM2_d
+ N_XXDEC/NET0141_XXDec/XI31/XI3/MM2_g N_VDD_XXDec/XI31/XI3/MM2_s
+ N_VDD_XXDec/XI31/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI30/XI3/MM2 N_XXDEC/XI30/XI3/NET13_XXDec/XI30/XI3/MM2_d
+ N_XXDEC/NET0141_XXDec/XI30/XI3/MM2_g N_VDD_XXDec/XI30/XI3/MM2_s
+ N_VDD_XXDec/XI30/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI27/XI3/MM2 N_XXDEC/XI27/XI3/NET13_XXDec/XI27/XI3/MM2_d
+ N_XXDEC/NET0141_XXDec/XI27/XI3/MM2_g N_VDD_XXDec/XI27/XI3/MM2_s
+ N_VDD_XXDec/XI27/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI36/XI3/MM3 N_WL<59>_XXDec/XI36/XI3/MM3_d
+ N_XXDEC/NET0123_XXDec/XI36/XI3/MM3_g
+ N_XXDEC/XI36/XI3/NET13_XXDec/XI36/XI3/MM3_s N_VDD_XXDec/XI36/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI3/MM3 N_WL<51>_XXDec/XI35/XI3/MM3_d
+ N_XXDEC/NET187_XXDec/XI35/XI3/MM3_g
+ N_XXDEC/XI35/XI3/NET13_XXDec/XI35/XI3/MM3_s N_VDD_XXDec/XI35/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI3/MM3 N_WL<43>_XXDec/XI34/XI3/MM3_d
+ N_XXDEC/NET188_XXDec/XI34/XI3/MM3_g
+ N_XXDEC/XI34/XI3/NET13_XXDec/XI34/XI3/MM3_s N_VDD_XXDec/XI34/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI3/MM3 N_WL<35>_XXDec/XI33/XI3/MM3_d
+ N_XXDEC/NET0122_XXDec/XI33/XI3/MM3_g
+ N_XXDEC/XI33/XI3/NET13_XXDec/XI33/XI3/MM3_s N_VDD_XXDec/XI33/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI3/MM3 N_WL<27>_XXDec/XI32/XI3/MM3_d
+ N_XXDEC/NET190_XXDec/XI32/XI3/MM3_g
+ N_XXDEC/XI32/XI3/NET13_XXDec/XI32/XI3/MM3_s N_VDD_XXDec/XI32/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI3/MM3 N_WL<19>_XXDec/XI31/XI3/MM3_d
+ N_XXDEC/NET0220_XXDec/XI31/XI3/MM3_g
+ N_XXDEC/XI31/XI3/NET13_XXDec/XI31/XI3/MM3_s N_VDD_XXDec/XI31/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI3/MM3 N_WL<11>_XXDec/XI30/XI3/MM3_d
+ N_XXDEC/NET192_XXDec/XI30/XI3/MM3_g
+ N_XXDEC/XI30/XI3/NET13_XXDec/XI30/XI3/MM3_s N_VDD_XXDec/XI30/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI3/MM3 N_WL<3>_XXDec/XI27/XI3/MM3_d
+ N_XXDEC/NET0130_XXDec/XI27/XI3/MM3_g
+ N_XXDEC/XI27/XI3/NET13_XXDec/XI27/XI3/MM3_s N_VDD_XXDec/XI27/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI2/MM2 N_XXDEC/XI36/XI2/NET13_XXDec/XI36/XI2/MM2_d
+ N_XXDEC/NET0142_XXDec/XI36/XI2/MM2_g N_VDD_XXDec/XI36/XI2/MM2_s
+ N_VDD_XXDec/XI36/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI35/XI2/MM2 N_XXDEC/XI35/XI2/NET13_XXDec/XI35/XI2/MM2_d
+ N_XXDEC/NET0142_XXDec/XI35/XI2/MM2_g N_VDD_XXDec/XI35/XI2/MM2_s
+ N_VDD_XXDec/XI35/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI34/XI2/MM2 N_XXDEC/XI34/XI2/NET13_XXDec/XI34/XI2/MM2_d
+ N_XXDEC/NET0142_XXDec/XI34/XI2/MM2_g N_VDD_XXDec/XI34/XI2/MM2_s
+ N_VDD_XXDec/XI34/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI33/XI2/MM2 N_XXDEC/XI33/XI2/NET13_XXDec/XI33/XI2/MM2_d
+ N_XXDEC/NET0142_XXDec/XI33/XI2/MM2_g N_VDD_XXDec/XI33/XI2/MM2_s
+ N_VDD_XXDec/XI33/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI32/XI2/MM2 N_XXDEC/XI32/XI2/NET13_XXDec/XI32/XI2/MM2_d
+ N_XXDEC/NET0142_XXDec/XI32/XI2/MM2_g N_VDD_XXDec/XI32/XI2/MM2_s
+ N_VDD_XXDec/XI32/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI31/XI2/MM2 N_XXDEC/XI31/XI2/NET13_XXDec/XI31/XI2/MM2_d
+ N_XXDEC/NET0142_XXDec/XI31/XI2/MM2_g N_VDD_XXDec/XI31/XI2/MM2_s
+ N_VDD_XXDec/XI31/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI30/XI2/MM2 N_XXDEC/XI30/XI2/NET13_XXDec/XI30/XI2/MM2_d
+ N_XXDEC/NET0142_XXDec/XI30/XI2/MM2_g N_VDD_XXDec/XI30/XI2/MM2_s
+ N_VDD_XXDec/XI30/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI27/XI2/MM2 N_XXDEC/XI27/XI2/NET13_XXDec/XI27/XI2/MM2_d
+ N_XXDEC/NET0142_XXDec/XI27/XI2/MM2_g N_VDD_XXDec/XI27/XI2/MM2_s
+ N_VDD_XXDec/XI27/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI36/XI2/MM3 N_WL<58>_XXDec/XI36/XI2/MM3_d
+ N_XXDEC/NET0123_XXDec/XI36/XI2/MM3_g
+ N_XXDEC/XI36/XI2/NET13_XXDec/XI36/XI2/MM3_s N_VDD_XXDec/XI36/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI2/MM3 N_WL<50>_XXDec/XI35/XI2/MM3_d
+ N_XXDEC/NET187_XXDec/XI35/XI2/MM3_g
+ N_XXDEC/XI35/XI2/NET13_XXDec/XI35/XI2/MM3_s N_VDD_XXDec/XI35/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI2/MM3 N_WL<42>_XXDec/XI34/XI2/MM3_d
+ N_XXDEC/NET188_XXDec/XI34/XI2/MM3_g
+ N_XXDEC/XI34/XI2/NET13_XXDec/XI34/XI2/MM3_s N_VDD_XXDec/XI34/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI2/MM3 N_WL<34>_XXDec/XI33/XI2/MM3_d
+ N_XXDEC/NET0122_XXDec/XI33/XI2/MM3_g
+ N_XXDEC/XI33/XI2/NET13_XXDec/XI33/XI2/MM3_s N_VDD_XXDec/XI33/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI2/MM3 N_WL<26>_XXDec/XI32/XI2/MM3_d
+ N_XXDEC/NET190_XXDec/XI32/XI2/MM3_g
+ N_XXDEC/XI32/XI2/NET13_XXDec/XI32/XI2/MM3_s N_VDD_XXDec/XI32/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI2/MM3 N_WL<18>_XXDec/XI31/XI2/MM3_d
+ N_XXDEC/NET0220_XXDec/XI31/XI2/MM3_g
+ N_XXDEC/XI31/XI2/NET13_XXDec/XI31/XI2/MM3_s N_VDD_XXDec/XI31/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI2/MM3 N_WL<10>_XXDec/XI30/XI2/MM3_d
+ N_XXDEC/NET192_XXDec/XI30/XI2/MM3_g
+ N_XXDEC/XI30/XI2/NET13_XXDec/XI30/XI2/MM3_s N_VDD_XXDec/XI30/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI2/MM3 N_WL<2>_XXDec/XI27/XI2/MM3_d
+ N_XXDEC/NET0130_XXDec/XI27/XI2/MM3_g
+ N_XXDEC/XI27/XI2/NET13_XXDec/XI27/XI2/MM3_s N_VDD_XXDec/XI27/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI1/MM2 N_XXDEC/XI36/XI1/NET13_XXDec/XI36/XI1/MM2_d
+ N_XXDEC/NET0143_XXDec/XI36/XI1/MM2_g N_VDD_XXDec/XI36/XI1/MM2_s
+ N_VDD_XXDec/XI36/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI35/XI1/MM2 N_XXDEC/XI35/XI1/NET13_XXDec/XI35/XI1/MM2_d
+ N_XXDEC/NET0143_XXDec/XI35/XI1/MM2_g N_VDD_XXDec/XI35/XI1/MM2_s
+ N_VDD_XXDec/XI35/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI34/XI1/MM2 N_XXDEC/XI34/XI1/NET13_XXDec/XI34/XI1/MM2_d
+ N_XXDEC/NET0143_XXDec/XI34/XI1/MM2_g N_VDD_XXDec/XI34/XI1/MM2_s
+ N_VDD_XXDec/XI34/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI33/XI1/MM2 N_XXDEC/XI33/XI1/NET13_XXDec/XI33/XI1/MM2_d
+ N_XXDEC/NET0143_XXDec/XI33/XI1/MM2_g N_VDD_XXDec/XI33/XI1/MM2_s
+ N_VDD_XXDec/XI33/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI32/XI1/MM2 N_XXDEC/XI32/XI1/NET13_XXDec/XI32/XI1/MM2_d
+ N_XXDEC/NET0143_XXDec/XI32/XI1/MM2_g N_VDD_XXDec/XI32/XI1/MM2_s
+ N_VDD_XXDec/XI32/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI31/XI1/MM2 N_XXDEC/XI31/XI1/NET13_XXDec/XI31/XI1/MM2_d
+ N_XXDEC/NET0143_XXDec/XI31/XI1/MM2_g N_VDD_XXDec/XI31/XI1/MM2_s
+ N_VDD_XXDec/XI31/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI30/XI1/MM2 N_XXDEC/XI30/XI1/NET13_XXDec/XI30/XI1/MM2_d
+ N_XXDEC/NET0143_XXDec/XI30/XI1/MM2_g N_VDD_XXDec/XI30/XI1/MM2_s
+ N_VDD_XXDec/XI30/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI27/XI1/MM2 N_XXDEC/XI27/XI1/NET13_XXDec/XI27/XI1/MM2_d
+ N_XXDEC/NET0143_XXDec/XI27/XI1/MM2_g N_VDD_XXDec/XI27/XI1/MM2_s
+ N_VDD_XXDec/XI27/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI36/XI1/MM3 N_WL<57>_XXDec/XI36/XI1/MM3_d
+ N_XXDEC/NET0123_XXDec/XI36/XI1/MM3_g
+ N_XXDEC/XI36/XI1/NET13_XXDec/XI36/XI1/MM3_s N_VDD_XXDec/XI36/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI1/MM3 N_WL<49>_XXDec/XI35/XI1/MM3_d
+ N_XXDEC/NET187_XXDec/XI35/XI1/MM3_g
+ N_XXDEC/XI35/XI1/NET13_XXDec/XI35/XI1/MM3_s N_VDD_XXDec/XI35/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI1/MM3 N_WL<41>_XXDec/XI34/XI1/MM3_d
+ N_XXDEC/NET188_XXDec/XI34/XI1/MM3_g
+ N_XXDEC/XI34/XI1/NET13_XXDec/XI34/XI1/MM3_s N_VDD_XXDec/XI34/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI1/MM3 N_WL<33>_XXDec/XI33/XI1/MM3_d
+ N_XXDEC/NET0122_XXDec/XI33/XI1/MM3_g
+ N_XXDEC/XI33/XI1/NET13_XXDec/XI33/XI1/MM3_s N_VDD_XXDec/XI33/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI1/MM3 N_WL<25>_XXDec/XI32/XI1/MM3_d
+ N_XXDEC/NET190_XXDec/XI32/XI1/MM3_g
+ N_XXDEC/XI32/XI1/NET13_XXDec/XI32/XI1/MM3_s N_VDD_XXDec/XI32/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI1/MM3 N_WL<17>_XXDec/XI31/XI1/MM3_d
+ N_XXDEC/NET0220_XXDec/XI31/XI1/MM3_g
+ N_XXDEC/XI31/XI1/NET13_XXDec/XI31/XI1/MM3_s N_VDD_XXDec/XI31/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI1/MM3 N_WL<9>_XXDec/XI30/XI1/MM3_d
+ N_XXDEC/NET192_XXDec/XI30/XI1/MM3_g
+ N_XXDEC/XI30/XI1/NET13_XXDec/XI30/XI1/MM3_s N_VDD_XXDec/XI30/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI1/MM3 N_WL<1>_XXDec/XI27/XI1/MM3_d
+ N_XXDEC/NET0130_XXDec/XI27/XI1/MM3_g
+ N_XXDEC/XI27/XI1/NET13_XXDec/XI27/XI1/MM3_s N_VDD_XXDec/XI27/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI36/XI0/MM2 N_XXDEC/XI36/XI0/NET13_XXDec/XI36/XI0/MM2_d
+ N_XXDEC/NET0144_XXDec/XI36/XI0/MM2_g N_VDD_XXDec/XI36/XI0/MM2_s
+ N_VDD_XXDec/XI36/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI35/XI0/MM2 N_XXDEC/XI35/XI0/NET13_XXDec/XI35/XI0/MM2_d
+ N_XXDEC/NET0144_XXDec/XI35/XI0/MM2_g N_VDD_XXDec/XI35/XI0/MM2_s
+ N_VDD_XXDec/XI35/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI34/XI0/MM2 N_XXDEC/XI34/XI0/NET13_XXDec/XI34/XI0/MM2_d
+ N_XXDEC/NET0144_XXDec/XI34/XI0/MM2_g N_VDD_XXDec/XI34/XI0/MM2_s
+ N_VDD_XXDec/XI34/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI33/XI0/MM2 N_XXDEC/XI33/XI0/NET13_XXDec/XI33/XI0/MM2_d
+ N_XXDEC/NET0144_XXDec/XI33/XI0/MM2_g N_VDD_XXDec/XI33/XI0/MM2_s
+ N_VDD_XXDec/XI33/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI32/XI0/MM2 N_XXDEC/XI32/XI0/NET13_XXDec/XI32/XI0/MM2_d
+ N_XXDEC/NET0144_XXDec/XI32/XI0/MM2_g N_VDD_XXDec/XI32/XI0/MM2_s
+ N_VDD_XXDec/XI32/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI31/XI0/MM2 N_XXDEC/XI31/XI0/NET13_XXDec/XI31/XI0/MM2_d
+ N_XXDEC/NET0144_XXDec/XI31/XI0/MM2_g N_VDD_XXDec/XI31/XI0/MM2_s
+ N_VDD_XXDec/XI31/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI30/XI0/MM2 N_XXDEC/XI30/XI0/NET13_XXDec/XI30/XI0/MM2_d
+ N_XXDEC/NET0144_XXDec/XI30/XI0/MM2_g N_VDD_XXDec/XI30/XI0/MM2_s
+ N_VDD_XXDec/XI30/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI27/XI0/MM2 N_XXDEC/XI27/XI0/NET13_XXDec/XI27/XI0/MM2_d
+ N_XXDEC/NET0144_XXDec/XI27/XI0/MM2_g N_VDD_XXDec/XI27/XI0/MM2_s
+ N_VDD_XXDec/XI27/XI7/MM2_b P_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13
+ PD=5.1e-07 PS=1.48e-06
mXXDec/XI36/XI0/MM3 N_WL<56>_XXDec/XI36/XI0/MM3_d
+ N_XXDEC/NET0123_XXDec/XI36/XI0/MM3_g
+ N_XXDEC/XI36/XI0/NET13_XXDec/XI36/XI0/MM3_s N_VDD_XXDec/XI36/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI35/XI0/MM3 N_WL<48>_XXDec/XI35/XI0/MM3_d
+ N_XXDEC/NET187_XXDec/XI35/XI0/MM3_g
+ N_XXDEC/XI35/XI0/NET13_XXDec/XI35/XI0/MM3_s N_VDD_XXDec/XI35/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI34/XI0/MM3 N_WL<40>_XXDec/XI34/XI0/MM3_d
+ N_XXDEC/NET188_XXDec/XI34/XI0/MM3_g
+ N_XXDEC/XI34/XI0/NET13_XXDec/XI34/XI0/MM3_s N_VDD_XXDec/XI34/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI33/XI0/MM3 N_WL<32>_XXDec/XI33/XI0/MM3_d
+ N_XXDEC/NET0122_XXDec/XI33/XI0/MM3_g
+ N_XXDEC/XI33/XI0/NET13_XXDec/XI33/XI0/MM3_s N_VDD_XXDec/XI33/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI32/XI0/MM3 N_WL<24>_XXDec/XI32/XI0/MM3_d
+ N_XXDEC/NET190_XXDec/XI32/XI0/MM3_g
+ N_XXDEC/XI32/XI0/NET13_XXDec/XI32/XI0/MM3_s N_VDD_XXDec/XI32/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI31/XI0/MM3 N_WL<16>_XXDec/XI31/XI0/MM3_d
+ N_XXDEC/NET0220_XXDec/XI31/XI0/MM3_g
+ N_XXDEC/XI31/XI0/NET13_XXDec/XI31/XI0/MM3_s N_VDD_XXDec/XI31/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI30/XI0/MM3 N_WL<8>_XXDec/XI30/XI0/MM3_d
+ N_XXDEC/NET192_XXDec/XI30/XI0/MM3_g
+ N_XXDEC/XI30/XI0/NET13_XXDec/XI30/XI0/MM3_s N_VDD_XXDec/XI30/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXXDec/XI27/XI0/MM3 N_WL<0>_XXDec/XI27/XI0/MM3_d
+ N_XXDEC/NET0130_XXDec/XI27/XI0/MM3_g
+ N_XXDEC/XI27/XI0/NET13_XXDec/XI27/XI0/MM3_s N_VDD_XXDec/XI27/XI7/MM2_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07
mXROM/XI7/XI3/MM8 N_BL<0>_XROM/XI7/XI3/MM8_d N_WL<63>_XROM/XI7/XI3/MM8_g
+ N_VSS_XROM/XI7/XI3/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM6 XROM/XI7/XI3/NET119 N_WL<62>_XROM/XI7/XI3/MM6_g
+ N_VSS_XROM/XI7/XI3/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM8 N_BL<0>_XROM/XI7/XI2/MM8_d N_WL<61>_XROM/XI7/XI2/MM8_g
+ N_VSS_XROM/XI7/XI2/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM0 XROM/XI7/XI2/NET143 N_WL<60>_XROM/XI7/XI2/MM0_g
+ N_VSS_XROM/XI7/XI2/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM8 N_BL<0>_XROM/XI7/XI1/MM8_d N_WL<59>_XROM/XI7/XI1/MM8_g
+ N_VSS_XROM/XI7/XI1/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM0 XROM/XI7/XI1/NET143 N_WL<58>_XROM/XI7/XI1/MM0_g
+ N_VSS_XROM/XI7/XI1/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM8 N_BL<0>_XROM/XI7/XI0/MM8_d N_WL<57>_XROM/XI7/XI0/MM8_g
+ N_VSS_XROM/XI7/XI0/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM0 XROM/XI7/XI0/NET143 N_WL<56>_XROM/XI7/XI0/MM0_g
+ N_VSS_XROM/XI7/XI0/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM8 N_BL<0>_XROM/XI6/XI3/MM8_d N_WL<55>_XROM/XI6/XI3/MM8_g
+ N_VSS_XROM/XI6/XI3/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM0 XROM/XI6/XI3/NET143 N_WL<54>_XROM/XI6/XI3/MM0_g
+ N_VSS_XROM/XI6/XI3/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM8 N_BL<0>_XROM/XI6/XI2/MM8_d N_WL<53>_XROM/XI6/XI2/MM8_g
+ N_VSS_XROM/XI6/XI2/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM0 XROM/XI6/XI2/NET143 N_WL<52>_XROM/XI6/XI2/MM0_g
+ N_VSS_XROM/XI6/XI2/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM8 N_BL<0>_XROM/XI6/XI1/MM8_d N_WL<51>_XROM/XI6/XI1/MM8_g
+ N_VSS_XROM/XI6/XI1/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM0 XROM/XI6/XI1/NET143 N_WL<50>_XROM/XI6/XI1/MM0_g
+ N_VSS_XROM/XI6/XI1/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM8 N_BL<0>_XROM/XI6/XI0/MM8_d N_WL<49>_XROM/XI6/XI0/MM8_g
+ N_VSS_XROM/XI6/XI0/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM0 XROM/XI6/XI0/NET143 N_WL<48>_XROM/XI6/XI0/MM0_g
+ N_VSS_XROM/XI6/XI0/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM9 XROM/XI7/XI3/NET107 N_WL<63>_XROM/XI7/XI3/MM9_g
+ N_VSS_XROM/XI7/XI3/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM1 N_BL<1>_XROM/XI7/XI3/MM1_d N_WL<62>_XROM/XI7/XI3/MM1_g
+ N_VSS_XROM/XI7/XI3/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM9 XROM/XI7/XI2/NET107 N_WL<61>_XROM/XI7/XI2/MM9_g
+ N_VSS_XROM/XI7/XI2/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM1 N_BL<1>_XROM/XI7/XI2/MM1_d N_WL<60>_XROM/XI7/XI2/MM1_g
+ N_VSS_XROM/XI7/XI2/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM9 XROM/XI7/XI1/NET107 N_WL<59>_XROM/XI7/XI1/MM9_g
+ N_VSS_XROM/XI7/XI1/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM1 N_BL<1>_XROM/XI7/XI1/MM1_d N_WL<58>_XROM/XI7/XI1/MM1_g
+ N_VSS_XROM/XI7/XI1/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM9 XROM/XI7/XI0/NET107 N_WL<57>_XROM/XI7/XI0/MM9_g
+ N_VSS_XROM/XI7/XI0/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM1 N_BL<1>_XROM/XI7/XI0/MM1_d N_WL<56>_XROM/XI7/XI0/MM1_g
+ N_VSS_XROM/XI7/XI0/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM9 XROM/XI6/XI3/NET107 N_WL<55>_XROM/XI6/XI3/MM9_g
+ N_VSS_XROM/XI6/XI3/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM1 N_BL<1>_XROM/XI6/XI3/MM1_d N_WL<54>_XROM/XI6/XI3/MM1_g
+ N_VSS_XROM/XI6/XI3/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM9 XROM/XI6/XI2/NET107 N_WL<53>_XROM/XI6/XI2/MM9_g
+ N_VSS_XROM/XI6/XI2/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM1 N_BL<1>_XROM/XI6/XI2/MM1_d N_WL<52>_XROM/XI6/XI2/MM1_g
+ N_VSS_XROM/XI6/XI2/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM9 XROM/XI6/XI1/NET107 N_WL<51>_XROM/XI6/XI1/MM9_g
+ N_VSS_XROM/XI6/XI1/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM1 N_BL<1>_XROM/XI6/XI1/MM1_d N_WL<50>_XROM/XI6/XI1/MM1_g
+ N_VSS_XROM/XI6/XI1/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM9 XROM/XI6/XI0/NET107 N_WL<49>_XROM/XI6/XI0/MM9_g
+ N_VSS_XROM/XI6/XI0/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM1 N_BL<1>_XROM/XI6/XI0/MM1_d N_WL<48>_XROM/XI6/XI0/MM1_g
+ N_VSS_XROM/XI6/XI0/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM10 N_BL<2>_XROM/XI7/XI3/MM10_d N_WL<63>_XROM/XI7/XI3/MM10_g
+ N_VSS_XROM/XI7/XI3/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM2 XROM/XI7/XI7/NET135 N_WL<62>_XROM/XI7/XI7/MM2_g
+ N_VSS_XROM/XI7/XI7/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM10 N_BL<2>_XROM/XI7/XI2/MM10_d N_WL<61>_XROM/XI7/XI2/MM10_g
+ N_VSS_XROM/XI7/XI2/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM2 XROM/XI7/XI2/NET135 N_WL<60>_XROM/XI7/XI2/MM2_g
+ N_VSS_XROM/XI7/XI2/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM10 N_BL<2>_XROM/XI7/XI1/MM10_d N_WL<59>_XROM/XI7/XI1/MM10_g
+ N_VSS_XROM/XI7/XI1/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM2 XROM/XI7/XI1/NET135 N_WL<58>_XROM/XI7/XI1/MM2_g
+ N_VSS_XROM/XI7/XI1/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM10 N_BL<2>_XROM/XI7/XI0/MM10_d N_WL<57>_XROM/XI7/XI0/MM10_g
+ N_VSS_XROM/XI7/XI0/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM2 XROM/XI7/XI0/NET135 N_WL<56>_XROM/XI7/XI0/MM2_g
+ N_VSS_XROM/XI7/XI0/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM10 N_BL<2>_XROM/XI6/XI3/MM10_d N_WL<55>_XROM/XI6/XI3/MM10_g
+ N_VSS_XROM/XI6/XI3/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM2 XROM/XI6/XI3/NET135 N_WL<54>_XROM/XI6/XI3/MM2_g
+ N_VSS_XROM/XI6/XI3/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM10 N_BL<2>_XROM/XI6/XI2/MM10_d N_WL<53>_XROM/XI6/XI2/MM10_g
+ N_VSS_XROM/XI6/XI2/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM2 XROM/XI6/XI2/NET135 N_WL<52>_XROM/XI6/XI2/MM2_g
+ N_VSS_XROM/XI6/XI2/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM10 N_BL<2>_XROM/XI6/XI1/MM10_d N_WL<51>_XROM/XI6/XI1/MM10_g
+ N_VSS_XROM/XI6/XI1/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM2 XROM/XI6/XI1/NET135 N_WL<50>_XROM/XI6/XI1/MM2_g
+ N_VSS_XROM/XI6/XI1/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM10 N_BL<2>_XROM/XI6/XI0/MM10_d N_WL<49>_XROM/XI6/XI0/MM10_g
+ N_VSS_XROM/XI6/XI0/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM2 XROM/XI6/XI0/NET135 N_WL<48>_XROM/XI6/XI0/MM2_g
+ N_VSS_XROM/XI6/XI0/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM11 XROM/XI7/XI3/NET99 N_WL<63>_XROM/XI7/XI3/MM11_g
+ N_VSS_XROM/XI7/XI3/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM3 N_BL<3>_XROM/XI7/XI3/MM3_d N_WL<62>_XROM/XI7/XI3/MM3_g
+ N_VSS_XROM/XI7/XI3/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM11 XROM/XI7/XI2/NET99 N_WL<61>_XROM/XI7/XI2/MM11_g
+ N_VSS_XROM/XI7/XI2/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM3 N_BL<3>_XROM/XI7/XI2/MM3_d N_WL<60>_XROM/XI7/XI2/MM3_g
+ N_VSS_XROM/XI7/XI2/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM11 XROM/XI7/XI1/NET99 N_WL<59>_XROM/XI7/XI1/MM11_g
+ N_VSS_XROM/XI7/XI1/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM3 N_BL<3>_XROM/XI7/XI1/MM3_d N_WL<58>_XROM/XI7/XI1/MM3_g
+ N_VSS_XROM/XI7/XI1/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM11 XROM/XI7/XI0/NET99 N_WL<57>_XROM/XI7/XI0/MM11_g
+ N_VSS_XROM/XI7/XI0/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM3 N_BL<3>_XROM/XI7/XI0/MM3_d N_WL<56>_XROM/XI7/XI0/MM3_g
+ N_VSS_XROM/XI7/XI0/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM11 XROM/XI6/XI3/NET99 N_WL<55>_XROM/XI6/XI3/MM11_g
+ N_VSS_XROM/XI6/XI3/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM3 N_BL<3>_XROM/XI6/XI3/MM3_d N_WL<54>_XROM/XI6/XI3/MM3_g
+ N_VSS_XROM/XI6/XI3/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM11 XROM/XI6/XI2/NET99 N_WL<53>_XROM/XI6/XI2/MM11_g
+ N_VSS_XROM/XI6/XI2/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM3 N_BL<3>_XROM/XI6/XI2/MM3_d N_WL<52>_XROM/XI6/XI2/MM3_g
+ N_VSS_XROM/XI6/XI2/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM11 XROM/XI6/XI1/NET99 N_WL<51>_XROM/XI6/XI1/MM11_g
+ N_VSS_XROM/XI6/XI1/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM3 N_BL<3>_XROM/XI6/XI1/MM3_d N_WL<50>_XROM/XI6/XI1/MM3_g
+ N_VSS_XROM/XI6/XI1/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM11 XROM/XI6/XI0/NET99 N_WL<49>_XROM/XI6/XI0/MM11_g
+ N_VSS_XROM/XI6/XI0/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM3 N_BL<3>_XROM/XI6/XI0/MM3_d N_WL<48>_XROM/XI6/XI0/MM3_g
+ N_VSS_XROM/XI6/XI0/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM12 N_BL<4>_XROM/XI7/XI3/MM12_d N_WL<63>_XROM/XI7/XI3/MM12_g
+ N_VSS_XROM/XI7/XI3/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM2 XROM/XI7/XI3/NET135 N_WL<62>_XROM/XI7/XI3/MM2_g
+ N_VSS_XROM/XI7/XI3/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM12 N_BL<4>_XROM/XI7/XI2/MM12_d N_WL<61>_XROM/XI7/XI2/MM12_g
+ N_VSS_XROM/XI7/XI2/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM4 XROM/XI7/XI2/NET127 N_WL<60>_XROM/XI7/XI2/MM4_g
+ N_VSS_XROM/XI7/XI2/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM12 N_BL<4>_XROM/XI7/XI1/MM12_d N_WL<59>_XROM/XI7/XI1/MM12_g
+ N_VSS_XROM/XI7/XI1/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM4 XROM/XI7/XI1/NET127 N_WL<58>_XROM/XI7/XI1/MM4_g
+ N_VSS_XROM/XI7/XI1/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM12 N_BL<4>_XROM/XI7/XI0/MM12_d N_WL<57>_XROM/XI7/XI0/MM12_g
+ N_VSS_XROM/XI7/XI0/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM4 XROM/XI7/XI0/NET127 N_WL<56>_XROM/XI7/XI0/MM4_g
+ N_VSS_XROM/XI7/XI0/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM12 N_BL<4>_XROM/XI6/XI3/MM12_d N_WL<55>_XROM/XI6/XI3/MM12_g
+ N_VSS_XROM/XI6/XI3/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM4 XROM/XI6/XI3/NET127 N_WL<54>_XROM/XI6/XI3/MM4_g
+ N_VSS_XROM/XI6/XI3/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM12 N_BL<4>_XROM/XI6/XI2/MM12_d N_WL<53>_XROM/XI6/XI2/MM12_g
+ N_VSS_XROM/XI6/XI2/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM4 XROM/XI6/XI2/NET127 N_WL<52>_XROM/XI6/XI2/MM4_g
+ N_VSS_XROM/XI6/XI2/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM12 N_BL<4>_XROM/XI6/XI1/MM12_d N_WL<51>_XROM/XI6/XI1/MM12_g
+ N_VSS_XROM/XI6/XI1/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM4 XROM/XI6/XI1/NET127 N_WL<50>_XROM/XI6/XI1/MM4_g
+ N_VSS_XROM/XI6/XI1/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM12 N_BL<4>_XROM/XI6/XI0/MM12_d N_WL<49>_XROM/XI6/XI0/MM12_g
+ N_VSS_XROM/XI6/XI0/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM4 XROM/XI6/XI0/NET127 N_WL<48>_XROM/XI6/XI0/MM4_g
+ N_VSS_XROM/XI6/XI0/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM13 XROM/XI7/XI3/NET91 N_WL<63>_XROM/XI7/XI3/MM13_g
+ N_VSS_XROM/XI7/XI3/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM5 N_BL<5>_XROM/XI7/XI3/MM5_d N_WL<62>_XROM/XI7/XI3/MM5_g
+ N_VSS_XROM/XI7/XI3/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM13 XROM/XI7/XI2/NET91 N_WL<61>_XROM/XI7/XI2/MM13_g
+ N_VSS_XROM/XI7/XI2/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM5 N_BL<5>_XROM/XI7/XI2/MM5_d N_WL<60>_XROM/XI7/XI2/MM5_g
+ N_VSS_XROM/XI7/XI2/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM13 XROM/XI7/XI1/NET91 N_WL<59>_XROM/XI7/XI1/MM13_g
+ N_VSS_XROM/XI7/XI1/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM5 N_BL<5>_XROM/XI7/XI1/MM5_d N_WL<58>_XROM/XI7/XI1/MM5_g
+ N_VSS_XROM/XI7/XI1/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM13 XROM/XI7/XI0/NET91 N_WL<57>_XROM/XI7/XI0/MM13_g
+ N_VSS_XROM/XI7/XI0/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM5 N_BL<5>_XROM/XI7/XI0/MM5_d N_WL<56>_XROM/XI7/XI0/MM5_g
+ N_VSS_XROM/XI7/XI0/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM13 XROM/XI6/XI3/NET91 N_WL<55>_XROM/XI6/XI3/MM13_g
+ N_VSS_XROM/XI6/XI3/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM5 N_BL<5>_XROM/XI6/XI3/MM5_d N_WL<54>_XROM/XI6/XI3/MM5_g
+ N_VSS_XROM/XI6/XI3/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM13 XROM/XI6/XI2/NET91 N_WL<53>_XROM/XI6/XI2/MM13_g
+ N_VSS_XROM/XI6/XI2/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM5 N_BL<5>_XROM/XI6/XI2/MM5_d N_WL<52>_XROM/XI6/XI2/MM5_g
+ N_VSS_XROM/XI6/XI2/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM13 XROM/XI6/XI1/NET91 N_WL<51>_XROM/XI6/XI1/MM13_g
+ N_VSS_XROM/XI6/XI1/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM5 N_BL<5>_XROM/XI6/XI1/MM5_d N_WL<50>_XROM/XI6/XI1/MM5_g
+ N_VSS_XROM/XI6/XI1/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM13 XROM/XI6/XI0/NET91 N_WL<49>_XROM/XI6/XI0/MM13_g
+ N_VSS_XROM/XI6/XI0/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM5 N_BL<5>_XROM/XI6/XI0/MM5_d N_WL<48>_XROM/XI6/XI0/MM5_g
+ N_VSS_XROM/XI6/XI0/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM14 N_BL<6>_XROM/XI7/XI3/MM14_d N_WL<63>_XROM/XI7/XI3/MM14_g
+ N_VSS_XROM/XI7/XI3/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM6 XROM/XI7/XI7/NET119 N_WL<62>_XROM/XI7/XI7/MM6_g
+ N_VSS_XROM/XI7/XI7/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM14 N_BL<6>_XROM/XI7/XI2/MM14_d N_WL<61>_XROM/XI7/XI2/MM14_g
+ N_VSS_XROM/XI7/XI2/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM6 XROM/XI7/XI2/NET119 N_WL<60>_XROM/XI7/XI2/MM6_g
+ N_VSS_XROM/XI7/XI2/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM14 N_BL<6>_XROM/XI7/XI1/MM14_d N_WL<59>_XROM/XI7/XI1/MM14_g
+ N_VSS_XROM/XI7/XI1/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM6 XROM/XI7/XI1/NET119 N_WL<58>_XROM/XI7/XI1/MM6_g
+ N_VSS_XROM/XI7/XI1/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM14 N_BL<6>_XROM/XI7/XI0/MM14_d N_WL<57>_XROM/XI7/XI0/MM14_g
+ N_VSS_XROM/XI7/XI0/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM6 XROM/XI7/XI0/NET119 N_WL<56>_XROM/XI7/XI0/MM6_g
+ N_VSS_XROM/XI7/XI0/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM14 N_BL<6>_XROM/XI6/XI3/MM14_d N_WL<55>_XROM/XI6/XI3/MM14_g
+ N_VSS_XROM/XI6/XI3/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM6 XROM/XI6/XI3/NET119 N_WL<54>_XROM/XI6/XI3/MM6_g
+ N_VSS_XROM/XI6/XI3/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM14 N_BL<6>_XROM/XI6/XI2/MM14_d N_WL<53>_XROM/XI6/XI2/MM14_g
+ N_VSS_XROM/XI6/XI2/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM6 XROM/XI6/XI2/NET119 N_WL<52>_XROM/XI6/XI2/MM6_g
+ N_VSS_XROM/XI6/XI2/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM14 N_BL<6>_XROM/XI6/XI1/MM14_d N_WL<51>_XROM/XI6/XI1/MM14_g
+ N_VSS_XROM/XI6/XI1/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM6 XROM/XI6/XI1/NET119 N_WL<50>_XROM/XI6/XI1/MM6_g
+ N_VSS_XROM/XI6/XI1/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM14 N_BL<6>_XROM/XI6/XI0/MM14_d N_WL<49>_XROM/XI6/XI0/MM14_g
+ N_VSS_XROM/XI6/XI0/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM6 XROM/XI6/XI0/NET119 N_WL<48>_XROM/XI6/XI0/MM6_g
+ N_VSS_XROM/XI6/XI0/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM15 XROM/XI7/XI3/NET83 N_WL<63>_XROM/XI7/XI3/MM15_g
+ N_VSS_XROM/XI7/XI3/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM7 N_BL<7>_XROM/XI7/XI3/MM7_d N_WL<62>_XROM/XI7/XI3/MM7_g
+ N_VSS_XROM/XI7/XI3/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM15 XROM/XI7/XI2/NET83 N_WL<61>_XROM/XI7/XI2/MM15_g
+ N_VSS_XROM/XI7/XI2/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI2/MM7 N_BL<7>_XROM/XI7/XI2/MM7_d N_WL<60>_XROM/XI7/XI2/MM7_g
+ N_VSS_XROM/XI7/XI2/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM15 XROM/XI7/XI1/NET83 N_WL<59>_XROM/XI7/XI1/MM15_g
+ N_VSS_XROM/XI7/XI1/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI1/MM7 N_BL<7>_XROM/XI7/XI1/MM7_d N_WL<58>_XROM/XI7/XI1/MM7_g
+ N_VSS_XROM/XI7/XI1/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM15 XROM/XI7/XI0/NET83 N_WL<57>_XROM/XI7/XI0/MM15_g
+ N_VSS_XROM/XI7/XI0/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI0/MM7 N_BL<7>_XROM/XI7/XI0/MM7_d N_WL<56>_XROM/XI7/XI0/MM7_g
+ N_VSS_XROM/XI7/XI0/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM15 XROM/XI6/XI3/NET83 N_WL<55>_XROM/XI6/XI3/MM15_g
+ N_VSS_XROM/XI6/XI3/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI3/MM7 N_BL<7>_XROM/XI6/XI3/MM7_d N_WL<54>_XROM/XI6/XI3/MM7_g
+ N_VSS_XROM/XI6/XI3/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM15 XROM/XI6/XI2/NET83 N_WL<53>_XROM/XI6/XI2/MM15_g
+ N_VSS_XROM/XI6/XI2/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI2/MM7 N_BL<7>_XROM/XI6/XI2/MM7_d N_WL<52>_XROM/XI6/XI2/MM7_g
+ N_VSS_XROM/XI6/XI2/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM15 XROM/XI6/XI1/NET83 N_WL<51>_XROM/XI6/XI1/MM15_g
+ N_VSS_XROM/XI6/XI1/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI1/MM7 N_BL<7>_XROM/XI6/XI1/MM7_d N_WL<50>_XROM/XI6/XI1/MM7_g
+ N_VSS_XROM/XI6/XI1/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM15 XROM/XI6/XI0/NET83 N_WL<49>_XROM/XI6/XI0/MM15_g
+ N_VSS_XROM/XI6/XI0/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI0/MM7 N_BL<7>_XROM/XI6/XI0/MM7_d N_WL<48>_XROM/XI6/XI0/MM7_g
+ N_VSS_XROM/XI6/XI0/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM8 N_BL<8>_XROM/XI7/XI7/MM8_d N_WL<63>_XROM/XI7/XI7/MM8_g
+ N_VSS_XROM/XI7/XI7/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM4 XROM/XI7/XI3/NET127 N_WL<62>_XROM/XI7/XI3/MM4_g
+ N_VSS_XROM/XI7/XI3/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM8 N_BL<8>_XROM/XI7/XI6/MM8_d N_WL<61>_XROM/XI7/XI6/MM8_g
+ N_VSS_XROM/XI7/XI6/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM0 XROM/XI7/XI6/NET143 N_WL<60>_XROM/XI7/XI6/MM0_g
+ N_VSS_XROM/XI7/XI6/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM8 N_BL<8>_XROM/XI7/XI5/MM8_d N_WL<59>_XROM/XI7/XI5/MM8_g
+ N_VSS_XROM/XI7/XI5/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM0 XROM/XI7/XI5/NET143 N_WL<58>_XROM/XI7/XI5/MM0_g
+ N_VSS_XROM/XI7/XI5/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM8 N_BL<8>_XROM/XI7/XI4/MM8_d N_WL<57>_XROM/XI7/XI4/MM8_g
+ N_VSS_XROM/XI7/XI4/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM0 XROM/XI7/XI4/NET143 N_WL<56>_XROM/XI7/XI4/MM0_g
+ N_VSS_XROM/XI7/XI4/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM8 N_BL<8>_XROM/XI6/XI7/MM8_d N_WL<55>_XROM/XI6/XI7/MM8_g
+ N_VSS_XROM/XI6/XI7/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM0 XROM/XI6/XI7/NET143 N_WL<54>_XROM/XI6/XI7/MM0_g
+ N_VSS_XROM/XI6/XI7/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM8 N_BL<8>_XROM/XI6/XI6/MM8_d N_WL<53>_XROM/XI6/XI6/MM8_g
+ N_VSS_XROM/XI6/XI6/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM0 XROM/XI6/XI6/NET143 N_WL<52>_XROM/XI6/XI6/MM0_g
+ N_VSS_XROM/XI6/XI6/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM8 N_BL<8>_XROM/XI6/XI5/MM8_d N_WL<51>_XROM/XI6/XI5/MM8_g
+ N_VSS_XROM/XI6/XI5/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM0 XROM/XI6/XI5/NET143 N_WL<50>_XROM/XI6/XI5/MM0_g
+ N_VSS_XROM/XI6/XI5/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM8 N_BL<8>_XROM/XI6/XI4/MM8_d N_WL<49>_XROM/XI6/XI4/MM8_g
+ N_VSS_XROM/XI6/XI4/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM0 XROM/XI6/XI4/NET143 N_WL<48>_XROM/XI6/XI4/MM0_g
+ N_VSS_XROM/XI6/XI4/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM9 XROM/XI7/XI7/NET107 N_WL<63>_XROM/XI7/XI7/MM9_g
+ N_VSS_XROM/XI7/XI7/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM1 N_BL<9>_XROM/XI7/XI7/MM1_d N_WL<62>_XROM/XI7/XI7/MM1_g
+ N_VSS_XROM/XI7/XI7/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM9 XROM/XI7/XI6/NET107 N_WL<61>_XROM/XI7/XI6/MM9_g
+ N_VSS_XROM/XI7/XI6/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM1 N_BL<9>_XROM/XI7/XI6/MM1_d N_WL<60>_XROM/XI7/XI6/MM1_g
+ N_VSS_XROM/XI7/XI6/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM9 XROM/XI7/XI5/NET107 N_WL<59>_XROM/XI7/XI5/MM9_g
+ N_VSS_XROM/XI7/XI5/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM1 N_BL<9>_XROM/XI7/XI5/MM1_d N_WL<58>_XROM/XI7/XI5/MM1_g
+ N_VSS_XROM/XI7/XI5/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM9 XROM/XI7/XI4/NET107 N_WL<57>_XROM/XI7/XI4/MM9_g
+ N_VSS_XROM/XI7/XI4/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM1 N_BL<9>_XROM/XI7/XI4/MM1_d N_WL<56>_XROM/XI7/XI4/MM1_g
+ N_VSS_XROM/XI7/XI4/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM9 XROM/XI6/XI7/NET107 N_WL<55>_XROM/XI6/XI7/MM9_g
+ N_VSS_XROM/XI6/XI7/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM1 N_BL<9>_XROM/XI6/XI7/MM1_d N_WL<54>_XROM/XI6/XI7/MM1_g
+ N_VSS_XROM/XI6/XI7/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM9 XROM/XI6/XI6/NET107 N_WL<53>_XROM/XI6/XI6/MM9_g
+ N_VSS_XROM/XI6/XI6/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM1 N_BL<9>_XROM/XI6/XI6/MM1_d N_WL<52>_XROM/XI6/XI6/MM1_g
+ N_VSS_XROM/XI6/XI6/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM9 XROM/XI6/XI5/NET107 N_WL<51>_XROM/XI6/XI5/MM9_g
+ N_VSS_XROM/XI6/XI5/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM1 N_BL<9>_XROM/XI6/XI5/MM1_d N_WL<50>_XROM/XI6/XI5/MM1_g
+ N_VSS_XROM/XI6/XI5/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM9 XROM/XI6/XI4/NET107 N_WL<49>_XROM/XI6/XI4/MM9_g
+ N_VSS_XROM/XI6/XI4/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM1 N_BL<9>_XROM/XI6/XI4/MM1_d N_WL<48>_XROM/XI6/XI4/MM1_g
+ N_VSS_XROM/XI6/XI4/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM10 N_BL<10>_XROM/XI7/XI7/MM10_d N_WL<63>_XROM/XI7/XI7/MM10_g
+ N_VSS_XROM/XI7/XI7/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM4 XROM/XI7/XI7/NET127 N_WL<62>_XROM/XI7/XI7/MM4_g
+ N_VSS_XROM/XI7/XI7/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM10 N_BL<10>_XROM/XI7/XI6/MM10_d N_WL<61>_XROM/XI7/XI6/MM10_g
+ N_VSS_XROM/XI7/XI6/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM2 XROM/XI7/XI6/NET135 N_WL<60>_XROM/XI7/XI6/MM2_g
+ N_VSS_XROM/XI7/XI6/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM10 N_BL<10>_XROM/XI7/XI5/MM10_d N_WL<59>_XROM/XI7/XI5/MM10_g
+ N_VSS_XROM/XI7/XI5/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM2 XROM/XI7/XI5/NET135 N_WL<58>_XROM/XI7/XI5/MM2_g
+ N_VSS_XROM/XI7/XI5/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM10 N_BL<10>_XROM/XI7/XI4/MM10_d N_WL<57>_XROM/XI7/XI4/MM10_g
+ N_VSS_XROM/XI7/XI4/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM2 XROM/XI7/XI4/NET135 N_WL<56>_XROM/XI7/XI4/MM2_g
+ N_VSS_XROM/XI7/XI4/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM10 N_BL<10>_XROM/XI6/XI7/MM10_d N_WL<55>_XROM/XI6/XI7/MM10_g
+ N_VSS_XROM/XI6/XI7/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM2 XROM/XI6/XI7/NET135 N_WL<54>_XROM/XI6/XI7/MM2_g
+ N_VSS_XROM/XI6/XI7/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM10 N_BL<10>_XROM/XI6/XI6/MM10_d N_WL<53>_XROM/XI6/XI6/MM10_g
+ N_VSS_XROM/XI6/XI6/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM2 XROM/XI6/XI6/NET135 N_WL<52>_XROM/XI6/XI6/MM2_g
+ N_VSS_XROM/XI6/XI6/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM10 N_BL<10>_XROM/XI6/XI5/MM10_d N_WL<51>_XROM/XI6/XI5/MM10_g
+ N_VSS_XROM/XI6/XI5/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM2 XROM/XI6/XI5/NET135 N_WL<50>_XROM/XI6/XI5/MM2_g
+ N_VSS_XROM/XI6/XI5/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM10 N_BL<10>_XROM/XI6/XI4/MM10_d N_WL<49>_XROM/XI6/XI4/MM10_g
+ N_VSS_XROM/XI6/XI4/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM2 XROM/XI6/XI4/NET135 N_WL<48>_XROM/XI6/XI4/MM2_g
+ N_VSS_XROM/XI6/XI4/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM11 XROM/XI7/XI7/NET99 N_WL<63>_XROM/XI7/XI7/MM11_g
+ N_VSS_XROM/XI7/XI7/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM3 N_BL<11>_XROM/XI7/XI7/MM3_d N_WL<62>_XROM/XI7/XI7/MM3_g
+ N_VSS_XROM/XI7/XI7/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM11 XROM/XI7/XI6/NET99 N_WL<61>_XROM/XI7/XI6/MM11_g
+ N_VSS_XROM/XI7/XI6/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM3 N_BL<11>_XROM/XI7/XI6/MM3_d N_WL<60>_XROM/XI7/XI6/MM3_g
+ N_VSS_XROM/XI7/XI6/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM11 XROM/XI7/XI5/NET99 N_WL<59>_XROM/XI7/XI5/MM11_g
+ N_VSS_XROM/XI7/XI5/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM3 N_BL<11>_XROM/XI7/XI5/MM3_d N_WL<58>_XROM/XI7/XI5/MM3_g
+ N_VSS_XROM/XI7/XI5/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM11 XROM/XI7/XI4/NET99 N_WL<57>_XROM/XI7/XI4/MM11_g
+ N_VSS_XROM/XI7/XI4/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM3 N_BL<11>_XROM/XI7/XI4/MM3_d N_WL<56>_XROM/XI7/XI4/MM3_g
+ N_VSS_XROM/XI7/XI4/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM11 XROM/XI6/XI7/NET99 N_WL<55>_XROM/XI6/XI7/MM11_g
+ N_VSS_XROM/XI6/XI7/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM3 N_BL<11>_XROM/XI6/XI7/MM3_d N_WL<54>_XROM/XI6/XI7/MM3_g
+ N_VSS_XROM/XI6/XI7/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM11 XROM/XI6/XI6/NET99 N_WL<53>_XROM/XI6/XI6/MM11_g
+ N_VSS_XROM/XI6/XI6/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM3 N_BL<11>_XROM/XI6/XI6/MM3_d N_WL<52>_XROM/XI6/XI6/MM3_g
+ N_VSS_XROM/XI6/XI6/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM11 XROM/XI6/XI5/NET99 N_WL<51>_XROM/XI6/XI5/MM11_g
+ N_VSS_XROM/XI6/XI5/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM3 N_BL<11>_XROM/XI6/XI5/MM3_d N_WL<50>_XROM/XI6/XI5/MM3_g
+ N_VSS_XROM/XI6/XI5/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM11 XROM/XI6/XI4/NET99 N_WL<49>_XROM/XI6/XI4/MM11_g
+ N_VSS_XROM/XI6/XI4/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM3 N_BL<11>_XROM/XI6/XI4/MM3_d N_WL<48>_XROM/XI6/XI4/MM3_g
+ N_VSS_XROM/XI6/XI4/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM12 N_BL<12>_XROM/XI7/XI7/MM12_d N_WL<63>_XROM/XI7/XI7/MM12_g
+ N_VSS_XROM/XI7/XI7/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM0 XROM/XI7/XI7/NET143 N_WL<62>_XROM/XI7/XI7/MM0_g
+ N_VSS_XROM/XI7/XI7/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM12 N_BL<12>_XROM/XI7/XI6/MM12_d N_WL<61>_XROM/XI7/XI6/MM12_g
+ N_VSS_XROM/XI7/XI6/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM4 XROM/XI7/XI6/NET127 N_WL<60>_XROM/XI7/XI6/MM4_g
+ N_VSS_XROM/XI7/XI6/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM12 N_BL<12>_XROM/XI7/XI5/MM12_d N_WL<59>_XROM/XI7/XI5/MM12_g
+ N_VSS_XROM/XI7/XI5/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM4 XROM/XI7/XI5/NET127 N_WL<58>_XROM/XI7/XI5/MM4_g
+ N_VSS_XROM/XI7/XI5/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM12 N_BL<12>_XROM/XI7/XI4/MM12_d N_WL<57>_XROM/XI7/XI4/MM12_g
+ N_VSS_XROM/XI7/XI4/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM4 XROM/XI7/XI4/NET127 N_WL<56>_XROM/XI7/XI4/MM4_g
+ N_VSS_XROM/XI7/XI4/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM12 N_BL<12>_XROM/XI6/XI7/MM12_d N_WL<55>_XROM/XI6/XI7/MM12_g
+ N_VSS_XROM/XI6/XI7/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM4 XROM/XI6/XI7/NET127 N_WL<54>_XROM/XI6/XI7/MM4_g
+ N_VSS_XROM/XI6/XI7/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM12 N_BL<12>_XROM/XI6/XI6/MM12_d N_WL<53>_XROM/XI6/XI6/MM12_g
+ N_VSS_XROM/XI6/XI6/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM4 XROM/XI6/XI6/NET127 N_WL<52>_XROM/XI6/XI6/MM4_g
+ N_VSS_XROM/XI6/XI6/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM12 N_BL<12>_XROM/XI6/XI5/MM12_d N_WL<51>_XROM/XI6/XI5/MM12_g
+ N_VSS_XROM/XI6/XI5/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM4 XROM/XI6/XI5/NET127 N_WL<50>_XROM/XI6/XI5/MM4_g
+ N_VSS_XROM/XI6/XI5/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM12 N_BL<12>_XROM/XI6/XI4/MM12_d N_WL<49>_XROM/XI6/XI4/MM12_g
+ N_VSS_XROM/XI6/XI4/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM4 XROM/XI6/XI4/NET127 N_WL<48>_XROM/XI6/XI4/MM4_g
+ N_VSS_XROM/XI6/XI4/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM13 XROM/XI7/XI7/NET91 N_WL<63>_XROM/XI7/XI7/MM13_g
+ N_VSS_XROM/XI7/XI7/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM5 N_BL<13>_XROM/XI7/XI7/MM5_d N_WL<62>_XROM/XI7/XI7/MM5_g
+ N_VSS_XROM/XI7/XI7/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM13 XROM/XI7/XI6/NET91 N_WL<61>_XROM/XI7/XI6/MM13_g
+ N_VSS_XROM/XI7/XI6/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM5 N_BL<13>_XROM/XI7/XI6/MM5_d N_WL<60>_XROM/XI7/XI6/MM5_g
+ N_VSS_XROM/XI7/XI6/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM13 XROM/XI7/XI5/NET91 N_WL<59>_XROM/XI7/XI5/MM13_g
+ N_VSS_XROM/XI7/XI5/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM5 N_BL<13>_XROM/XI7/XI5/MM5_d N_WL<58>_XROM/XI7/XI5/MM5_g
+ N_VSS_XROM/XI7/XI5/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM13 XROM/XI7/XI4/NET91 N_WL<57>_XROM/XI7/XI4/MM13_g
+ N_VSS_XROM/XI7/XI4/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM5 N_BL<13>_XROM/XI7/XI4/MM5_d N_WL<56>_XROM/XI7/XI4/MM5_g
+ N_VSS_XROM/XI7/XI4/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM13 XROM/XI6/XI7/NET91 N_WL<55>_XROM/XI6/XI7/MM13_g
+ N_VSS_XROM/XI6/XI7/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM5 N_BL<13>_XROM/XI6/XI7/MM5_d N_WL<54>_XROM/XI6/XI7/MM5_g
+ N_VSS_XROM/XI6/XI7/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM13 XROM/XI6/XI6/NET91 N_WL<53>_XROM/XI6/XI6/MM13_g
+ N_VSS_XROM/XI6/XI6/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM5 N_BL<13>_XROM/XI6/XI6/MM5_d N_WL<52>_XROM/XI6/XI6/MM5_g
+ N_VSS_XROM/XI6/XI6/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM13 XROM/XI6/XI5/NET91 N_WL<51>_XROM/XI6/XI5/MM13_g
+ N_VSS_XROM/XI6/XI5/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM5 N_BL<13>_XROM/XI6/XI5/MM5_d N_WL<50>_XROM/XI6/XI5/MM5_g
+ N_VSS_XROM/XI6/XI5/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM13 XROM/XI6/XI4/NET91 N_WL<49>_XROM/XI6/XI4/MM13_g
+ N_VSS_XROM/XI6/XI4/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM5 N_BL<13>_XROM/XI6/XI4/MM5_d N_WL<48>_XROM/XI6/XI4/MM5_g
+ N_VSS_XROM/XI6/XI4/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM14 N_BL<14>_XROM/XI7/XI7/MM14_d N_WL<63>_XROM/XI7/XI7/MM14_g
+ N_VSS_XROM/XI7/XI7/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI3/MM0 XROM/XI7/XI3/NET143 N_WL<62>_XROM/XI7/XI3/MM0_g
+ N_VSS_XROM/XI7/XI3/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM14 N_BL<14>_XROM/XI7/XI6/MM14_d N_WL<61>_XROM/XI7/XI6/MM14_g
+ N_VSS_XROM/XI7/XI6/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM6 XROM/XI7/XI6/NET119 N_WL<60>_XROM/XI7/XI6/MM6_g
+ N_VSS_XROM/XI7/XI6/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM14 N_BL<14>_XROM/XI7/XI5/MM14_d N_WL<59>_XROM/XI7/XI5/MM14_g
+ N_VSS_XROM/XI7/XI5/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM6 XROM/XI7/XI5/NET119 N_WL<58>_XROM/XI7/XI5/MM6_g
+ N_VSS_XROM/XI7/XI5/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM14 N_BL<14>_XROM/XI7/XI4/MM14_d N_WL<57>_XROM/XI7/XI4/MM14_g
+ N_VSS_XROM/XI7/XI4/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM6 XROM/XI7/XI4/NET119 N_WL<56>_XROM/XI7/XI4/MM6_g
+ N_VSS_XROM/XI7/XI4/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM14 N_BL<14>_XROM/XI6/XI7/MM14_d N_WL<55>_XROM/XI6/XI7/MM14_g
+ N_VSS_XROM/XI6/XI7/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM6 XROM/XI6/XI7/NET119 N_WL<54>_XROM/XI6/XI7/MM6_g
+ N_VSS_XROM/XI6/XI7/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM14 N_BL<14>_XROM/XI6/XI6/MM14_d N_WL<53>_XROM/XI6/XI6/MM14_g
+ N_VSS_XROM/XI6/XI6/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM6 XROM/XI6/XI6/NET119 N_WL<52>_XROM/XI6/XI6/MM6_g
+ N_VSS_XROM/XI6/XI6/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM14 N_BL<14>_XROM/XI6/XI5/MM14_d N_WL<51>_XROM/XI6/XI5/MM14_g
+ N_VSS_XROM/XI6/XI5/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM6 XROM/XI6/XI5/NET119 N_WL<50>_XROM/XI6/XI5/MM6_g
+ N_VSS_XROM/XI6/XI5/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM14 N_BL<14>_XROM/XI6/XI4/MM14_d N_WL<49>_XROM/XI6/XI4/MM14_g
+ N_VSS_XROM/XI6/XI4/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM6 XROM/XI6/XI4/NET119 N_WL<48>_XROM/XI6/XI4/MM6_g
+ N_VSS_XROM/XI6/XI4/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM15 XROM/XI7/XI7/NET83 N_WL<63>_XROM/XI7/XI7/MM15_g
+ N_VSS_XROM/XI7/XI7/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI7/MM7 N_BL<15>_XROM/XI7/XI7/MM7_d N_WL<62>_XROM/XI7/XI7/MM7_g
+ N_VSS_XROM/XI7/XI7/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM15 XROM/XI7/XI6/NET83 N_WL<61>_XROM/XI7/XI6/MM15_g
+ N_VSS_XROM/XI7/XI6/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI6/MM7 N_BL<15>_XROM/XI7/XI6/MM7_d N_WL<60>_XROM/XI7/XI6/MM7_g
+ N_VSS_XROM/XI7/XI6/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM15 XROM/XI7/XI5/NET83 N_WL<59>_XROM/XI7/XI5/MM15_g
+ N_VSS_XROM/XI7/XI5/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI5/MM7 N_BL<15>_XROM/XI7/XI5/MM7_d N_WL<58>_XROM/XI7/XI5/MM7_g
+ N_VSS_XROM/XI7/XI5/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM15 XROM/XI7/XI4/NET83 N_WL<57>_XROM/XI7/XI4/MM15_g
+ N_VSS_XROM/XI7/XI4/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI7/XI4/MM7 N_BL<15>_XROM/XI7/XI4/MM7_d N_WL<56>_XROM/XI7/XI4/MM7_g
+ N_VSS_XROM/XI7/XI4/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM15 XROM/XI6/XI7/NET83 N_WL<55>_XROM/XI6/XI7/MM15_g
+ N_VSS_XROM/XI6/XI7/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI7/MM7 N_BL<15>_XROM/XI6/XI7/MM7_d N_WL<54>_XROM/XI6/XI7/MM7_g
+ N_VSS_XROM/XI6/XI7/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM15 XROM/XI6/XI6/NET83 N_WL<53>_XROM/XI6/XI6/MM15_g
+ N_VSS_XROM/XI6/XI6/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI6/MM7 N_BL<15>_XROM/XI6/XI6/MM7_d N_WL<52>_XROM/XI6/XI6/MM7_g
+ N_VSS_XROM/XI6/XI6/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM15 XROM/XI6/XI5/NET83 N_WL<51>_XROM/XI6/XI5/MM15_g
+ N_VSS_XROM/XI6/XI5/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI5/MM7 N_BL<15>_XROM/XI6/XI5/MM7_d N_WL<50>_XROM/XI6/XI5/MM7_g
+ N_VSS_XROM/XI6/XI5/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM15 XROM/XI6/XI4/NET83 N_WL<49>_XROM/XI6/XI4/MM15_g
+ N_VSS_XROM/XI6/XI4/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI6/XI4/MM7 N_BL<15>_XROM/XI6/XI4/MM7_d N_WL<48>_XROM/XI6/XI4/MM7_g
+ N_VSS_XROM/XI6/XI4/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM8 N_BL<0>_XROM/XI5/XI3/MM8_d N_WL<47>_XROM/XI5/XI3/MM8_g
+ N_VSS_XROM/XI5/XI3/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM0 XROM/XI5/XI3/NET143 N_WL<46>_XROM/XI5/XI3/MM0_g
+ N_VSS_XROM/XI5/XI3/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM8 N_BL<0>_XROM/XI5/XI2/MM8_d N_WL<45>_XROM/XI5/XI2/MM8_g
+ N_VSS_XROM/XI5/XI2/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM0 XROM/XI5/XI2/NET143 N_WL<44>_XROM/XI5/XI2/MM0_g
+ N_VSS_XROM/XI5/XI2/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM8 N_BL<0>_XROM/XI5/XI1/MM8_d N_WL<43>_XROM/XI5/XI1/MM8_g
+ N_VSS_XROM/XI5/XI1/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM0 XROM/XI5/XI1/NET143 N_WL<42>_XROM/XI5/XI1/MM0_g
+ N_VSS_XROM/XI5/XI1/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM8 N_BL<0>_XROM/XI5/XI0/MM8_d N_WL<41>_XROM/XI5/XI0/MM8_g
+ N_VSS_XROM/XI5/XI0/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM0 XROM/XI5/XI0/NET143 N_WL<40>_XROM/XI5/XI0/MM0_g
+ N_VSS_XROM/XI5/XI0/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM8 N_BL<0>_XROM/XI4/XI3/MM8_d N_WL<39>_XROM/XI4/XI3/MM8_g
+ N_VSS_XROM/XI4/XI3/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM0 XROM/XI4/XI3/NET143 N_WL<38>_XROM/XI4/XI3/MM0_g
+ N_VSS_XROM/XI4/XI3/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM8 N_BL<0>_XROM/XI4/XI2/MM8_d N_WL<37>_XROM/XI4/XI2/MM8_g
+ N_VSS_XROM/XI4/XI2/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM0 XROM/XI4/XI2/NET143 N_WL<36>_XROM/XI4/XI2/MM0_g
+ N_VSS_XROM/XI4/XI2/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM8 N_BL<0>_XROM/XI4/XI1/MM8_d N_WL<35>_XROM/XI4/XI1/MM8_g
+ N_VSS_XROM/XI4/XI1/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM0 XROM/XI4/XI1/NET143 N_WL<34>_XROM/XI4/XI1/MM0_g
+ N_VSS_XROM/XI4/XI1/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM8 N_BL<0>_XROM/XI4/XI0/MM8_d N_WL<33>_XROM/XI4/XI0/MM8_g
+ N_VSS_XROM/XI4/XI0/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM0 XROM/XI4/XI0/NET143 N_WL<32>_XROM/XI4/XI0/MM0_g
+ N_VSS_XROM/XI4/XI0/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM9 XROM/XI5/XI3/NET107 N_WL<47>_XROM/XI5/XI3/MM9_g
+ N_VSS_XROM/XI5/XI3/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM1 N_BL<1>_XROM/XI5/XI3/MM1_d N_WL<46>_XROM/XI5/XI3/MM1_g
+ N_VSS_XROM/XI5/XI3/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM9 XROM/XI5/XI2/NET107 N_WL<45>_XROM/XI5/XI2/MM9_g
+ N_VSS_XROM/XI5/XI2/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM1 N_BL<1>_XROM/XI5/XI2/MM1_d N_WL<44>_XROM/XI5/XI2/MM1_g
+ N_VSS_XROM/XI5/XI2/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM9 XROM/XI5/XI1/NET107 N_WL<43>_XROM/XI5/XI1/MM9_g
+ N_VSS_XROM/XI5/XI1/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM1 N_BL<1>_XROM/XI5/XI1/MM1_d N_WL<42>_XROM/XI5/XI1/MM1_g
+ N_VSS_XROM/XI5/XI1/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM9 XROM/XI5/XI0/NET107 N_WL<41>_XROM/XI5/XI0/MM9_g
+ N_VSS_XROM/XI5/XI0/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM1 N_BL<1>_XROM/XI5/XI0/MM1_d N_WL<40>_XROM/XI5/XI0/MM1_g
+ N_VSS_XROM/XI5/XI0/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM9 XROM/XI4/XI3/NET107 N_WL<39>_XROM/XI4/XI3/MM9_g
+ N_VSS_XROM/XI4/XI3/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM1 N_BL<1>_XROM/XI4/XI3/MM1_d N_WL<38>_XROM/XI4/XI3/MM1_g
+ N_VSS_XROM/XI4/XI3/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM9 XROM/XI4/XI2/NET107 N_WL<37>_XROM/XI4/XI2/MM9_g
+ N_VSS_XROM/XI4/XI2/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM1 N_BL<1>_XROM/XI4/XI2/MM1_d N_WL<36>_XROM/XI4/XI2/MM1_g
+ N_VSS_XROM/XI4/XI2/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM9 XROM/XI4/XI1/NET107 N_WL<35>_XROM/XI4/XI1/MM9_g
+ N_VSS_XROM/XI4/XI1/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM1 N_BL<1>_XROM/XI4/XI1/MM1_d N_WL<34>_XROM/XI4/XI1/MM1_g
+ N_VSS_XROM/XI4/XI1/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM9 XROM/XI4/XI0/NET107 N_WL<33>_XROM/XI4/XI0/MM9_g
+ N_VSS_XROM/XI4/XI0/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM1 N_BL<1>_XROM/XI4/XI0/MM1_d N_WL<32>_XROM/XI4/XI0/MM1_g
+ N_VSS_XROM/XI4/XI0/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM10 N_BL<2>_XROM/XI5/XI3/MM10_d N_WL<47>_XROM/XI5/XI3/MM10_g
+ N_VSS_XROM/XI5/XI3/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM2 XROM/XI5/XI3/NET135 N_WL<46>_XROM/XI5/XI3/MM2_g
+ N_VSS_XROM/XI5/XI3/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM10 N_BL<2>_XROM/XI5/XI2/MM10_d N_WL<45>_XROM/XI5/XI2/MM10_g
+ N_VSS_XROM/XI5/XI2/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM2 XROM/XI5/XI2/NET135 N_WL<44>_XROM/XI5/XI2/MM2_g
+ N_VSS_XROM/XI5/XI2/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM10 N_BL<2>_XROM/XI5/XI1/MM10_d N_WL<43>_XROM/XI5/XI1/MM10_g
+ N_VSS_XROM/XI5/XI1/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM2 XROM/XI5/XI1/NET135 N_WL<42>_XROM/XI5/XI1/MM2_g
+ N_VSS_XROM/XI5/XI1/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM10 N_BL<2>_XROM/XI5/XI0/MM10_d N_WL<41>_XROM/XI5/XI0/MM10_g
+ N_VSS_XROM/XI5/XI0/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM2 XROM/XI5/XI0/NET135 N_WL<40>_XROM/XI5/XI0/MM2_g
+ N_VSS_XROM/XI5/XI0/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM10 N_BL<2>_XROM/XI4/XI3/MM10_d N_WL<39>_XROM/XI4/XI3/MM10_g
+ N_VSS_XROM/XI4/XI3/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM2 XROM/XI4/XI3/NET135 N_WL<38>_XROM/XI4/XI3/MM2_g
+ N_VSS_XROM/XI4/XI3/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM10 N_BL<2>_XROM/XI4/XI2/MM10_d N_WL<37>_XROM/XI4/XI2/MM10_g
+ N_VSS_XROM/XI4/XI2/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM2 XROM/XI4/XI2/NET135 N_WL<36>_XROM/XI4/XI2/MM2_g
+ N_VSS_XROM/XI4/XI2/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM10 N_BL<2>_XROM/XI4/XI1/MM10_d N_WL<35>_XROM/XI4/XI1/MM10_g
+ N_VSS_XROM/XI4/XI1/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM2 XROM/XI4/XI1/NET135 N_WL<34>_XROM/XI4/XI1/MM2_g
+ N_VSS_XROM/XI4/XI1/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM10 N_BL<2>_XROM/XI4/XI0/MM10_d N_WL<33>_XROM/XI4/XI0/MM10_g
+ N_VSS_XROM/XI4/XI0/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM2 XROM/XI4/XI0/NET135 N_WL<32>_XROM/XI4/XI0/MM2_g
+ N_VSS_XROM/XI4/XI0/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM11 XROM/XI5/XI3/NET99 N_WL<47>_XROM/XI5/XI3/MM11_g
+ N_VSS_XROM/XI5/XI3/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM3 N_BL<3>_XROM/XI5/XI3/MM3_d N_WL<46>_XROM/XI5/XI3/MM3_g
+ N_VSS_XROM/XI5/XI3/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM11 XROM/XI5/XI2/NET99 N_WL<45>_XROM/XI5/XI2/MM11_g
+ N_VSS_XROM/XI5/XI2/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM3 N_BL<3>_XROM/XI5/XI2/MM3_d N_WL<44>_XROM/XI5/XI2/MM3_g
+ N_VSS_XROM/XI5/XI2/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM11 XROM/XI5/XI1/NET99 N_WL<43>_XROM/XI5/XI1/MM11_g
+ N_VSS_XROM/XI5/XI1/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM3 N_BL<3>_XROM/XI5/XI1/MM3_d N_WL<42>_XROM/XI5/XI1/MM3_g
+ N_VSS_XROM/XI5/XI1/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM11 XROM/XI5/XI0/NET99 N_WL<41>_XROM/XI5/XI0/MM11_g
+ N_VSS_XROM/XI5/XI0/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM3 N_BL<3>_XROM/XI5/XI0/MM3_d N_WL<40>_XROM/XI5/XI0/MM3_g
+ N_VSS_XROM/XI5/XI0/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM11 XROM/XI4/XI3/NET99 N_WL<39>_XROM/XI4/XI3/MM11_g
+ N_VSS_XROM/XI4/XI3/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM3 N_BL<3>_XROM/XI4/XI3/MM3_d N_WL<38>_XROM/XI4/XI3/MM3_g
+ N_VSS_XROM/XI4/XI3/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM11 XROM/XI4/XI2/NET99 N_WL<37>_XROM/XI4/XI2/MM11_g
+ N_VSS_XROM/XI4/XI2/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM3 N_BL<3>_XROM/XI4/XI2/MM3_d N_WL<36>_XROM/XI4/XI2/MM3_g
+ N_VSS_XROM/XI4/XI2/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM11 XROM/XI4/XI1/NET99 N_WL<35>_XROM/XI4/XI1/MM11_g
+ N_VSS_XROM/XI4/XI1/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM3 N_BL<3>_XROM/XI4/XI1/MM3_d N_WL<34>_XROM/XI4/XI1/MM3_g
+ N_VSS_XROM/XI4/XI1/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM11 XROM/XI4/XI0/NET99 N_WL<33>_XROM/XI4/XI0/MM11_g
+ N_VSS_XROM/XI4/XI0/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM3 N_BL<3>_XROM/XI4/XI0/MM3_d N_WL<32>_XROM/XI4/XI0/MM3_g
+ N_VSS_XROM/XI4/XI0/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM12 N_BL<4>_XROM/XI5/XI3/MM12_d N_WL<47>_XROM/XI5/XI3/MM12_g
+ N_VSS_XROM/XI5/XI3/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM4 XROM/XI5/XI3/NET127 N_WL<46>_XROM/XI5/XI3/MM4_g
+ N_VSS_XROM/XI5/XI3/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM12 N_BL<4>_XROM/XI5/XI2/MM12_d N_WL<45>_XROM/XI5/XI2/MM12_g
+ N_VSS_XROM/XI5/XI2/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM4 XROM/XI5/XI2/NET127 N_WL<44>_XROM/XI5/XI2/MM4_g
+ N_VSS_XROM/XI5/XI2/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM12 N_BL<4>_XROM/XI5/XI1/MM12_d N_WL<43>_XROM/XI5/XI1/MM12_g
+ N_VSS_XROM/XI5/XI1/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM4 XROM/XI5/XI1/NET127 N_WL<42>_XROM/XI5/XI1/MM4_g
+ N_VSS_XROM/XI5/XI1/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM12 N_BL<4>_XROM/XI5/XI0/MM12_d N_WL<41>_XROM/XI5/XI0/MM12_g
+ N_VSS_XROM/XI5/XI0/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM4 XROM/XI5/XI0/NET127 N_WL<40>_XROM/XI5/XI0/MM4_g
+ N_VSS_XROM/XI5/XI0/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM12 N_BL<4>_XROM/XI4/XI3/MM12_d N_WL<39>_XROM/XI4/XI3/MM12_g
+ N_VSS_XROM/XI4/XI3/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM4 XROM/XI4/XI3/NET127 N_WL<38>_XROM/XI4/XI3/MM4_g
+ N_VSS_XROM/XI4/XI3/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM12 N_BL<4>_XROM/XI4/XI2/MM12_d N_WL<37>_XROM/XI4/XI2/MM12_g
+ N_VSS_XROM/XI4/XI2/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM4 XROM/XI4/XI2/NET127 N_WL<36>_XROM/XI4/XI2/MM4_g
+ N_VSS_XROM/XI4/XI2/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM12 N_BL<4>_XROM/XI4/XI1/MM12_d N_WL<35>_XROM/XI4/XI1/MM12_g
+ N_VSS_XROM/XI4/XI1/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM4 XROM/XI4/XI1/NET127 N_WL<34>_XROM/XI4/XI1/MM4_g
+ N_VSS_XROM/XI4/XI1/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM12 N_BL<4>_XROM/XI4/XI0/MM12_d N_WL<33>_XROM/XI4/XI0/MM12_g
+ N_VSS_XROM/XI4/XI0/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM4 XROM/XI4/XI0/NET127 N_WL<32>_XROM/XI4/XI0/MM4_g
+ N_VSS_XROM/XI4/XI0/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM13 XROM/XI5/XI3/NET91 N_WL<47>_XROM/XI5/XI3/MM13_g
+ N_VSS_XROM/XI5/XI3/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM5 N_BL<5>_XROM/XI5/XI3/MM5_d N_WL<46>_XROM/XI5/XI3/MM5_g
+ N_VSS_XROM/XI5/XI3/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM13 XROM/XI5/XI2/NET91 N_WL<45>_XROM/XI5/XI2/MM13_g
+ N_VSS_XROM/XI5/XI2/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM5 N_BL<5>_XROM/XI5/XI2/MM5_d N_WL<44>_XROM/XI5/XI2/MM5_g
+ N_VSS_XROM/XI5/XI2/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM13 XROM/XI5/XI1/NET91 N_WL<43>_XROM/XI5/XI1/MM13_g
+ N_VSS_XROM/XI5/XI1/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM5 N_BL<5>_XROM/XI5/XI1/MM5_d N_WL<42>_XROM/XI5/XI1/MM5_g
+ N_VSS_XROM/XI5/XI1/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM13 XROM/XI5/XI0/NET91 N_WL<41>_XROM/XI5/XI0/MM13_g
+ N_VSS_XROM/XI5/XI0/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM5 N_BL<5>_XROM/XI5/XI0/MM5_d N_WL<40>_XROM/XI5/XI0/MM5_g
+ N_VSS_XROM/XI5/XI0/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM13 XROM/XI4/XI3/NET91 N_WL<39>_XROM/XI4/XI3/MM13_g
+ N_VSS_XROM/XI4/XI3/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM5 N_BL<5>_XROM/XI4/XI3/MM5_d N_WL<38>_XROM/XI4/XI3/MM5_g
+ N_VSS_XROM/XI4/XI3/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM13 XROM/XI4/XI2/NET91 N_WL<37>_XROM/XI4/XI2/MM13_g
+ N_VSS_XROM/XI4/XI2/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM5 N_BL<5>_XROM/XI4/XI2/MM5_d N_WL<36>_XROM/XI4/XI2/MM5_g
+ N_VSS_XROM/XI4/XI2/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM13 XROM/XI4/XI1/NET91 N_WL<35>_XROM/XI4/XI1/MM13_g
+ N_VSS_XROM/XI4/XI1/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM5 N_BL<5>_XROM/XI4/XI1/MM5_d N_WL<34>_XROM/XI4/XI1/MM5_g
+ N_VSS_XROM/XI4/XI1/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM13 XROM/XI4/XI0/NET91 N_WL<33>_XROM/XI4/XI0/MM13_g
+ N_VSS_XROM/XI4/XI0/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM5 N_BL<5>_XROM/XI4/XI0/MM5_d N_WL<32>_XROM/XI4/XI0/MM5_g
+ N_VSS_XROM/XI4/XI0/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM14 N_BL<6>_XROM/XI5/XI3/MM14_d N_WL<47>_XROM/XI5/XI3/MM14_g
+ N_VSS_XROM/XI5/XI3/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM6 XROM/XI5/XI3/NET119 N_WL<46>_XROM/XI5/XI3/MM6_g
+ N_VSS_XROM/XI5/XI3/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM14 N_BL<6>_XROM/XI5/XI2/MM14_d N_WL<45>_XROM/XI5/XI2/MM14_g
+ N_VSS_XROM/XI5/XI2/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM6 XROM/XI5/XI2/NET119 N_WL<44>_XROM/XI5/XI2/MM6_g
+ N_VSS_XROM/XI5/XI2/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM14 N_BL<6>_XROM/XI5/XI1/MM14_d N_WL<43>_XROM/XI5/XI1/MM14_g
+ N_VSS_XROM/XI5/XI1/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM6 XROM/XI5/XI1/NET119 N_WL<42>_XROM/XI5/XI1/MM6_g
+ N_VSS_XROM/XI5/XI1/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM14 N_BL<6>_XROM/XI5/XI0/MM14_d N_WL<41>_XROM/XI5/XI0/MM14_g
+ N_VSS_XROM/XI5/XI0/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM6 XROM/XI5/XI0/NET119 N_WL<40>_XROM/XI5/XI0/MM6_g
+ N_VSS_XROM/XI5/XI0/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM14 N_BL<6>_XROM/XI4/XI3/MM14_d N_WL<39>_XROM/XI4/XI3/MM14_g
+ N_VSS_XROM/XI4/XI3/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM6 XROM/XI4/XI3/NET119 N_WL<38>_XROM/XI4/XI3/MM6_g
+ N_VSS_XROM/XI4/XI3/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM14 N_BL<6>_XROM/XI4/XI2/MM14_d N_WL<37>_XROM/XI4/XI2/MM14_g
+ N_VSS_XROM/XI4/XI2/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM6 XROM/XI4/XI2/NET119 N_WL<36>_XROM/XI4/XI2/MM6_g
+ N_VSS_XROM/XI4/XI2/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM14 N_BL<6>_XROM/XI4/XI1/MM14_d N_WL<35>_XROM/XI4/XI1/MM14_g
+ N_VSS_XROM/XI4/XI1/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM6 XROM/XI4/XI1/NET119 N_WL<34>_XROM/XI4/XI1/MM6_g
+ N_VSS_XROM/XI4/XI1/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM14 N_BL<6>_XROM/XI4/XI0/MM14_d N_WL<33>_XROM/XI4/XI0/MM14_g
+ N_VSS_XROM/XI4/XI0/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM6 XROM/XI4/XI0/NET119 N_WL<32>_XROM/XI4/XI0/MM6_g
+ N_VSS_XROM/XI4/XI0/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM15 XROM/XI5/XI3/NET83 N_WL<47>_XROM/XI5/XI3/MM15_g
+ N_VSS_XROM/XI5/XI3/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI3/MM7 N_BL<7>_XROM/XI5/XI3/MM7_d N_WL<46>_XROM/XI5/XI3/MM7_g
+ N_VSS_XROM/XI5/XI3/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM15 XROM/XI5/XI2/NET83 N_WL<45>_XROM/XI5/XI2/MM15_g
+ N_VSS_XROM/XI5/XI2/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI2/MM7 N_BL<7>_XROM/XI5/XI2/MM7_d N_WL<44>_XROM/XI5/XI2/MM7_g
+ N_VSS_XROM/XI5/XI2/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM15 XROM/XI5/XI1/NET83 N_WL<43>_XROM/XI5/XI1/MM15_g
+ N_VSS_XROM/XI5/XI1/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI1/MM7 N_BL<7>_XROM/XI5/XI1/MM7_d N_WL<42>_XROM/XI5/XI1/MM7_g
+ N_VSS_XROM/XI5/XI1/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM15 XROM/XI5/XI0/NET83 N_WL<41>_XROM/XI5/XI0/MM15_g
+ N_VSS_XROM/XI5/XI0/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI0/MM7 N_BL<7>_XROM/XI5/XI0/MM7_d N_WL<40>_XROM/XI5/XI0/MM7_g
+ N_VSS_XROM/XI5/XI0/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM15 XROM/XI4/XI3/NET83 N_WL<39>_XROM/XI4/XI3/MM15_g
+ N_VSS_XROM/XI4/XI3/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI3/MM7 N_BL<7>_XROM/XI4/XI3/MM7_d N_WL<38>_XROM/XI4/XI3/MM7_g
+ N_VSS_XROM/XI4/XI3/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM15 XROM/XI4/XI2/NET83 N_WL<37>_XROM/XI4/XI2/MM15_g
+ N_VSS_XROM/XI4/XI2/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI2/MM7 N_BL<7>_XROM/XI4/XI2/MM7_d N_WL<36>_XROM/XI4/XI2/MM7_g
+ N_VSS_XROM/XI4/XI2/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM15 XROM/XI4/XI1/NET83 N_WL<35>_XROM/XI4/XI1/MM15_g
+ N_VSS_XROM/XI4/XI1/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI1/MM7 N_BL<7>_XROM/XI4/XI1/MM7_d N_WL<34>_XROM/XI4/XI1/MM7_g
+ N_VSS_XROM/XI4/XI1/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM15 XROM/XI4/XI0/NET83 N_WL<33>_XROM/XI4/XI0/MM15_g
+ N_VSS_XROM/XI4/XI0/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI0/MM7 N_BL<7>_XROM/XI4/XI0/MM7_d N_WL<32>_XROM/XI4/XI0/MM7_g
+ N_VSS_XROM/XI4/XI0/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM8 N_BL<8>_XROM/XI5/XI7/MM8_d N_WL<47>_XROM/XI5/XI7/MM8_g
+ N_VSS_XROM/XI5/XI7/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM0 XROM/XI5/XI7/NET143 N_WL<46>_XROM/XI5/XI7/MM0_g
+ N_VSS_XROM/XI5/XI7/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM8 N_BL<8>_XROM/XI5/XI6/MM8_d N_WL<45>_XROM/XI5/XI6/MM8_g
+ N_VSS_XROM/XI5/XI6/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM0 XROM/XI5/XI6/NET143 N_WL<44>_XROM/XI5/XI6/MM0_g
+ N_VSS_XROM/XI5/XI6/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM8 N_BL<8>_XROM/XI5/XI5/MM8_d N_WL<43>_XROM/XI5/XI5/MM8_g
+ N_VSS_XROM/XI5/XI5/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM0 XROM/XI5/XI5/NET143 N_WL<42>_XROM/XI5/XI5/MM0_g
+ N_VSS_XROM/XI5/XI5/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM8 N_BL<8>_XROM/XI5/XI4/MM8_d N_WL<41>_XROM/XI5/XI4/MM8_g
+ N_VSS_XROM/XI5/XI4/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM0 XROM/XI5/XI4/NET143 N_WL<40>_XROM/XI5/XI4/MM0_g
+ N_VSS_XROM/XI5/XI4/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM8 N_BL<8>_XROM/XI4/XI7/MM8_d N_WL<39>_XROM/XI4/XI7/MM8_g
+ N_VSS_XROM/XI4/XI7/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM0 XROM/XI4/XI7/NET143 N_WL<38>_XROM/XI4/XI7/MM0_g
+ N_VSS_XROM/XI4/XI7/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM8 N_BL<8>_XROM/XI4/XI6/MM8_d N_WL<37>_XROM/XI4/XI6/MM8_g
+ N_VSS_XROM/XI4/XI6/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM0 XROM/XI4/XI6/NET143 N_WL<36>_XROM/XI4/XI6/MM0_g
+ N_VSS_XROM/XI4/XI6/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM8 N_BL<8>_XROM/XI4/XI5/MM8_d N_WL<35>_XROM/XI4/XI5/MM8_g
+ N_VSS_XROM/XI4/XI5/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM0 XROM/XI4/XI5/NET143 N_WL<34>_XROM/XI4/XI5/MM0_g
+ N_VSS_XROM/XI4/XI5/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM8 N_BL<8>_XROM/XI4/XI4/MM8_d N_WL<33>_XROM/XI4/XI4/MM8_g
+ N_VSS_XROM/XI4/XI4/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM0 XROM/XI4/XI4/NET143 N_WL<32>_XROM/XI4/XI4/MM0_g
+ N_VSS_XROM/XI4/XI4/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM9 XROM/XI5/XI7/NET107 N_WL<47>_XROM/XI5/XI7/MM9_g
+ N_VSS_XROM/XI5/XI7/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM1 N_BL<9>_XROM/XI5/XI7/MM1_d N_WL<46>_XROM/XI5/XI7/MM1_g
+ N_VSS_XROM/XI5/XI7/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM9 XROM/XI5/XI6/NET107 N_WL<45>_XROM/XI5/XI6/MM9_g
+ N_VSS_XROM/XI5/XI6/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM1 N_BL<9>_XROM/XI5/XI6/MM1_d N_WL<44>_XROM/XI5/XI6/MM1_g
+ N_VSS_XROM/XI5/XI6/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM9 XROM/XI5/XI5/NET107 N_WL<43>_XROM/XI5/XI5/MM9_g
+ N_VSS_XROM/XI5/XI5/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM1 N_BL<9>_XROM/XI5/XI5/MM1_d N_WL<42>_XROM/XI5/XI5/MM1_g
+ N_VSS_XROM/XI5/XI5/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM9 XROM/XI5/XI4/NET107 N_WL<41>_XROM/XI5/XI4/MM9_g
+ N_VSS_XROM/XI5/XI4/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM1 N_BL<9>_XROM/XI5/XI4/MM1_d N_WL<40>_XROM/XI5/XI4/MM1_g
+ N_VSS_XROM/XI5/XI4/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM9 XROM/XI4/XI7/NET107 N_WL<39>_XROM/XI4/XI7/MM9_g
+ N_VSS_XROM/XI4/XI7/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM1 N_BL<9>_XROM/XI4/XI7/MM1_d N_WL<38>_XROM/XI4/XI7/MM1_g
+ N_VSS_XROM/XI4/XI7/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM9 XROM/XI4/XI6/NET107 N_WL<37>_XROM/XI4/XI6/MM9_g
+ N_VSS_XROM/XI4/XI6/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM1 N_BL<9>_XROM/XI4/XI6/MM1_d N_WL<36>_XROM/XI4/XI6/MM1_g
+ N_VSS_XROM/XI4/XI6/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM9 XROM/XI4/XI5/NET107 N_WL<35>_XROM/XI4/XI5/MM9_g
+ N_VSS_XROM/XI4/XI5/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM1 N_BL<9>_XROM/XI4/XI5/MM1_d N_WL<34>_XROM/XI4/XI5/MM1_g
+ N_VSS_XROM/XI4/XI5/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM9 XROM/XI4/XI4/NET107 N_WL<33>_XROM/XI4/XI4/MM9_g
+ N_VSS_XROM/XI4/XI4/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM1 N_BL<9>_XROM/XI4/XI4/MM1_d N_WL<32>_XROM/XI4/XI4/MM1_g
+ N_VSS_XROM/XI4/XI4/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM10 N_BL<10>_XROM/XI5/XI7/MM10_d N_WL<47>_XROM/XI5/XI7/MM10_g
+ N_VSS_XROM/XI5/XI7/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM2 XROM/XI5/XI7/NET135 N_WL<46>_XROM/XI5/XI7/MM2_g
+ N_VSS_XROM/XI5/XI7/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM10 N_BL<10>_XROM/XI5/XI6/MM10_d N_WL<45>_XROM/XI5/XI6/MM10_g
+ N_VSS_XROM/XI5/XI6/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM2 XROM/XI5/XI6/NET135 N_WL<44>_XROM/XI5/XI6/MM2_g
+ N_VSS_XROM/XI5/XI6/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM10 N_BL<10>_XROM/XI5/XI5/MM10_d N_WL<43>_XROM/XI5/XI5/MM10_g
+ N_VSS_XROM/XI5/XI5/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM2 XROM/XI5/XI5/NET135 N_WL<42>_XROM/XI5/XI5/MM2_g
+ N_VSS_XROM/XI5/XI5/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM10 N_BL<10>_XROM/XI5/XI4/MM10_d N_WL<41>_XROM/XI5/XI4/MM10_g
+ N_VSS_XROM/XI5/XI4/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM2 XROM/XI5/XI4/NET135 N_WL<40>_XROM/XI5/XI4/MM2_g
+ N_VSS_XROM/XI5/XI4/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM10 N_BL<10>_XROM/XI4/XI7/MM10_d N_WL<39>_XROM/XI4/XI7/MM10_g
+ N_VSS_XROM/XI4/XI7/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM2 XROM/XI4/XI7/NET135 N_WL<38>_XROM/XI4/XI7/MM2_g
+ N_VSS_XROM/XI4/XI7/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM10 N_BL<10>_XROM/XI4/XI6/MM10_d N_WL<37>_XROM/XI4/XI6/MM10_g
+ N_VSS_XROM/XI4/XI6/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM2 XROM/XI4/XI6/NET135 N_WL<36>_XROM/XI4/XI6/MM2_g
+ N_VSS_XROM/XI4/XI6/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM10 N_BL<10>_XROM/XI4/XI5/MM10_d N_WL<35>_XROM/XI4/XI5/MM10_g
+ N_VSS_XROM/XI4/XI5/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM2 XROM/XI4/XI5/NET135 N_WL<34>_XROM/XI4/XI5/MM2_g
+ N_VSS_XROM/XI4/XI5/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM10 N_BL<10>_XROM/XI4/XI4/MM10_d N_WL<33>_XROM/XI4/XI4/MM10_g
+ N_VSS_XROM/XI4/XI4/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM2 XROM/XI4/XI4/NET135 N_WL<32>_XROM/XI4/XI4/MM2_g
+ N_VSS_XROM/XI4/XI4/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM11 XROM/XI5/XI7/NET99 N_WL<47>_XROM/XI5/XI7/MM11_g
+ N_VSS_XROM/XI5/XI7/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM3 N_BL<11>_XROM/XI5/XI7/MM3_d N_WL<46>_XROM/XI5/XI7/MM3_g
+ N_VSS_XROM/XI5/XI7/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM11 XROM/XI5/XI6/NET99 N_WL<45>_XROM/XI5/XI6/MM11_g
+ N_VSS_XROM/XI5/XI6/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM3 N_BL<11>_XROM/XI5/XI6/MM3_d N_WL<44>_XROM/XI5/XI6/MM3_g
+ N_VSS_XROM/XI5/XI6/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM11 XROM/XI5/XI5/NET99 N_WL<43>_XROM/XI5/XI5/MM11_g
+ N_VSS_XROM/XI5/XI5/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM3 N_BL<11>_XROM/XI5/XI5/MM3_d N_WL<42>_XROM/XI5/XI5/MM3_g
+ N_VSS_XROM/XI5/XI5/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM11 XROM/XI5/XI4/NET99 N_WL<41>_XROM/XI5/XI4/MM11_g
+ N_VSS_XROM/XI5/XI4/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM3 N_BL<11>_XROM/XI5/XI4/MM3_d N_WL<40>_XROM/XI5/XI4/MM3_g
+ N_VSS_XROM/XI5/XI4/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM11 XROM/XI4/XI7/NET99 N_WL<39>_XROM/XI4/XI7/MM11_g
+ N_VSS_XROM/XI4/XI7/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM3 N_BL<11>_XROM/XI4/XI7/MM3_d N_WL<38>_XROM/XI4/XI7/MM3_g
+ N_VSS_XROM/XI4/XI7/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM11 XROM/XI4/XI6/NET99 N_WL<37>_XROM/XI4/XI6/MM11_g
+ N_VSS_XROM/XI4/XI6/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM3 N_BL<11>_XROM/XI4/XI6/MM3_d N_WL<36>_XROM/XI4/XI6/MM3_g
+ N_VSS_XROM/XI4/XI6/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM11 XROM/XI4/XI5/NET99 N_WL<35>_XROM/XI4/XI5/MM11_g
+ N_VSS_XROM/XI4/XI5/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM3 N_BL<11>_XROM/XI4/XI5/MM3_d N_WL<34>_XROM/XI4/XI5/MM3_g
+ N_VSS_XROM/XI4/XI5/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM11 XROM/XI4/XI4/NET99 N_WL<33>_XROM/XI4/XI4/MM11_g
+ N_VSS_XROM/XI4/XI4/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM3 N_BL<11>_XROM/XI4/XI4/MM3_d N_WL<32>_XROM/XI4/XI4/MM3_g
+ N_VSS_XROM/XI4/XI4/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM12 N_BL<12>_XROM/XI5/XI7/MM12_d N_WL<47>_XROM/XI5/XI7/MM12_g
+ N_VSS_XROM/XI5/XI7/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM4 XROM/XI5/XI7/NET127 N_WL<46>_XROM/XI5/XI7/MM4_g
+ N_VSS_XROM/XI5/XI7/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM12 N_BL<12>_XROM/XI5/XI6/MM12_d N_WL<45>_XROM/XI5/XI6/MM12_g
+ N_VSS_XROM/XI5/XI6/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM4 XROM/XI5/XI6/NET127 N_WL<44>_XROM/XI5/XI6/MM4_g
+ N_VSS_XROM/XI5/XI6/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM12 N_BL<12>_XROM/XI5/XI5/MM12_d N_WL<43>_XROM/XI5/XI5/MM12_g
+ N_VSS_XROM/XI5/XI5/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM4 XROM/XI5/XI5/NET127 N_WL<42>_XROM/XI5/XI5/MM4_g
+ N_VSS_XROM/XI5/XI5/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM12 N_BL<12>_XROM/XI5/XI4/MM12_d N_WL<41>_XROM/XI5/XI4/MM12_g
+ N_VSS_XROM/XI5/XI4/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM4 XROM/XI5/XI4/NET127 N_WL<40>_XROM/XI5/XI4/MM4_g
+ N_VSS_XROM/XI5/XI4/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM12 N_BL<12>_XROM/XI4/XI7/MM12_d N_WL<39>_XROM/XI4/XI7/MM12_g
+ N_VSS_XROM/XI4/XI7/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM4 XROM/XI4/XI7/NET127 N_WL<38>_XROM/XI4/XI7/MM4_g
+ N_VSS_XROM/XI4/XI7/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM12 N_BL<12>_XROM/XI4/XI6/MM12_d N_WL<37>_XROM/XI4/XI6/MM12_g
+ N_VSS_XROM/XI4/XI6/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM4 XROM/XI4/XI6/NET127 N_WL<36>_XROM/XI4/XI6/MM4_g
+ N_VSS_XROM/XI4/XI6/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM12 N_BL<12>_XROM/XI4/XI5/MM12_d N_WL<35>_XROM/XI4/XI5/MM12_g
+ N_VSS_XROM/XI4/XI5/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM4 XROM/XI4/XI5/NET127 N_WL<34>_XROM/XI4/XI5/MM4_g
+ N_VSS_XROM/XI4/XI5/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM12 N_BL<12>_XROM/XI4/XI4/MM12_d N_WL<33>_XROM/XI4/XI4/MM12_g
+ N_VSS_XROM/XI4/XI4/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM4 XROM/XI4/XI4/NET127 N_WL<32>_XROM/XI4/XI4/MM4_g
+ N_VSS_XROM/XI4/XI4/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM13 XROM/XI5/XI7/NET91 N_WL<47>_XROM/XI5/XI7/MM13_g
+ N_VSS_XROM/XI5/XI7/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM5 N_BL<13>_XROM/XI5/XI7/MM5_d N_WL<46>_XROM/XI5/XI7/MM5_g
+ N_VSS_XROM/XI5/XI7/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM13 XROM/XI5/XI6/NET91 N_WL<45>_XROM/XI5/XI6/MM13_g
+ N_VSS_XROM/XI5/XI6/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM5 N_BL<13>_XROM/XI5/XI6/MM5_d N_WL<44>_XROM/XI5/XI6/MM5_g
+ N_VSS_XROM/XI5/XI6/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM13 XROM/XI5/XI5/NET91 N_WL<43>_XROM/XI5/XI5/MM13_g
+ N_VSS_XROM/XI5/XI5/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM5 N_BL<13>_XROM/XI5/XI5/MM5_d N_WL<42>_XROM/XI5/XI5/MM5_g
+ N_VSS_XROM/XI5/XI5/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM13 XROM/XI5/XI4/NET91 N_WL<41>_XROM/XI5/XI4/MM13_g
+ N_VSS_XROM/XI5/XI4/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM5 N_BL<13>_XROM/XI5/XI4/MM5_d N_WL<40>_XROM/XI5/XI4/MM5_g
+ N_VSS_XROM/XI5/XI4/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM13 XROM/XI4/XI7/NET91 N_WL<39>_XROM/XI4/XI7/MM13_g
+ N_VSS_XROM/XI4/XI7/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM5 N_BL<13>_XROM/XI4/XI7/MM5_d N_WL<38>_XROM/XI4/XI7/MM5_g
+ N_VSS_XROM/XI4/XI7/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM13 XROM/XI4/XI6/NET91 N_WL<37>_XROM/XI4/XI6/MM13_g
+ N_VSS_XROM/XI4/XI6/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM5 N_BL<13>_XROM/XI4/XI6/MM5_d N_WL<36>_XROM/XI4/XI6/MM5_g
+ N_VSS_XROM/XI4/XI6/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM13 XROM/XI4/XI5/NET91 N_WL<35>_XROM/XI4/XI5/MM13_g
+ N_VSS_XROM/XI4/XI5/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM5 N_BL<13>_XROM/XI4/XI5/MM5_d N_WL<34>_XROM/XI4/XI5/MM5_g
+ N_VSS_XROM/XI4/XI5/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM13 XROM/XI4/XI4/NET91 N_WL<33>_XROM/XI4/XI4/MM13_g
+ N_VSS_XROM/XI4/XI4/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM5 N_BL<13>_XROM/XI4/XI4/MM5_d N_WL<32>_XROM/XI4/XI4/MM5_g
+ N_VSS_XROM/XI4/XI4/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM14 N_BL<14>_XROM/XI5/XI7/MM14_d N_WL<47>_XROM/XI5/XI7/MM14_g
+ N_VSS_XROM/XI5/XI7/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM6 XROM/XI5/XI7/NET119 N_WL<46>_XROM/XI5/XI7/MM6_g
+ N_VSS_XROM/XI5/XI7/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM14 N_BL<14>_XROM/XI5/XI6/MM14_d N_WL<45>_XROM/XI5/XI6/MM14_g
+ N_VSS_XROM/XI5/XI6/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM6 XROM/XI5/XI6/NET119 N_WL<44>_XROM/XI5/XI6/MM6_g
+ N_VSS_XROM/XI5/XI6/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM14 N_BL<14>_XROM/XI5/XI5/MM14_d N_WL<43>_XROM/XI5/XI5/MM14_g
+ N_VSS_XROM/XI5/XI5/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM6 XROM/XI5/XI5/NET119 N_WL<42>_XROM/XI5/XI5/MM6_g
+ N_VSS_XROM/XI5/XI5/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM14 N_BL<14>_XROM/XI5/XI4/MM14_d N_WL<41>_XROM/XI5/XI4/MM14_g
+ N_VSS_XROM/XI5/XI4/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM6 XROM/XI5/XI4/NET119 N_WL<40>_XROM/XI5/XI4/MM6_g
+ N_VSS_XROM/XI5/XI4/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM14 N_BL<14>_XROM/XI4/XI7/MM14_d N_WL<39>_XROM/XI4/XI7/MM14_g
+ N_VSS_XROM/XI4/XI7/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM6 XROM/XI4/XI7/NET119 N_WL<38>_XROM/XI4/XI7/MM6_g
+ N_VSS_XROM/XI4/XI7/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM14 N_BL<14>_XROM/XI4/XI6/MM14_d N_WL<37>_XROM/XI4/XI6/MM14_g
+ N_VSS_XROM/XI4/XI6/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM6 XROM/XI4/XI6/NET119 N_WL<36>_XROM/XI4/XI6/MM6_g
+ N_VSS_XROM/XI4/XI6/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM14 N_BL<14>_XROM/XI4/XI5/MM14_d N_WL<35>_XROM/XI4/XI5/MM14_g
+ N_VSS_XROM/XI4/XI5/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM6 XROM/XI4/XI5/NET119 N_WL<34>_XROM/XI4/XI5/MM6_g
+ N_VSS_XROM/XI4/XI5/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM14 N_BL<14>_XROM/XI4/XI4/MM14_d N_WL<33>_XROM/XI4/XI4/MM14_g
+ N_VSS_XROM/XI4/XI4/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM6 XROM/XI4/XI4/NET119 N_WL<32>_XROM/XI4/XI4/MM6_g
+ N_VSS_XROM/XI4/XI4/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM15 XROM/XI5/XI7/NET83 N_WL<47>_XROM/XI5/XI7/MM15_g
+ N_VSS_XROM/XI5/XI7/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI7/MM7 N_BL<15>_XROM/XI5/XI7/MM7_d N_WL<46>_XROM/XI5/XI7/MM7_g
+ N_VSS_XROM/XI5/XI7/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM15 XROM/XI5/XI6/NET83 N_WL<45>_XROM/XI5/XI6/MM15_g
+ N_VSS_XROM/XI5/XI6/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI6/MM7 N_BL<15>_XROM/XI5/XI6/MM7_d N_WL<44>_XROM/XI5/XI6/MM7_g
+ N_VSS_XROM/XI5/XI6/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM15 XROM/XI5/XI5/NET83 N_WL<43>_XROM/XI5/XI5/MM15_g
+ N_VSS_XROM/XI5/XI5/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI5/MM7 N_BL<15>_XROM/XI5/XI5/MM7_d N_WL<42>_XROM/XI5/XI5/MM7_g
+ N_VSS_XROM/XI5/XI5/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM15 XROM/XI5/XI4/NET83 N_WL<41>_XROM/XI5/XI4/MM15_g
+ N_VSS_XROM/XI5/XI4/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI5/XI4/MM7 N_BL<15>_XROM/XI5/XI4/MM7_d N_WL<40>_XROM/XI5/XI4/MM7_g
+ N_VSS_XROM/XI5/XI4/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM15 XROM/XI4/XI7/NET83 N_WL<39>_XROM/XI4/XI7/MM15_g
+ N_VSS_XROM/XI4/XI7/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI7/MM7 N_BL<15>_XROM/XI4/XI7/MM7_d N_WL<38>_XROM/XI4/XI7/MM7_g
+ N_VSS_XROM/XI4/XI7/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM15 XROM/XI4/XI6/NET83 N_WL<37>_XROM/XI4/XI6/MM15_g
+ N_VSS_XROM/XI4/XI6/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI6/MM7 N_BL<15>_XROM/XI4/XI6/MM7_d N_WL<36>_XROM/XI4/XI6/MM7_g
+ N_VSS_XROM/XI4/XI6/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM15 XROM/XI4/XI5/NET83 N_WL<35>_XROM/XI4/XI5/MM15_g
+ N_VSS_XROM/XI4/XI5/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI5/MM7 N_BL<15>_XROM/XI4/XI5/MM7_d N_WL<34>_XROM/XI4/XI5/MM7_g
+ N_VSS_XROM/XI4/XI5/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM15 XROM/XI4/XI4/NET83 N_WL<33>_XROM/XI4/XI4/MM15_g
+ N_VSS_XROM/XI4/XI4/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI4/XI4/MM7 N_BL<15>_XROM/XI4/XI4/MM7_d N_WL<32>_XROM/XI4/XI4/MM7_g
+ N_VSS_XROM/XI4/XI4/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM8 N_BL<0>_XROM/XI3/XI3/MM8_d N_WL<31>_XROM/XI3/XI3/MM8_g
+ N_VSS_XROM/XI3/XI3/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM0 XROM/XI3/XI3/NET143 N_WL<30>_XROM/XI3/XI3/MM0_g
+ N_VSS_XROM/XI3/XI3/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM8 N_BL<0>_XROM/XI3/XI2/MM8_d N_WL<29>_XROM/XI3/XI2/MM8_g
+ N_VSS_XROM/XI3/XI2/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM0 XROM/XI3/XI2/NET143 N_WL<28>_XROM/XI3/XI2/MM0_g
+ N_VSS_XROM/XI3/XI2/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM8 N_BL<0>_XROM/XI3/XI1/MM8_d N_WL<27>_XROM/XI3/XI1/MM8_g
+ N_VSS_XROM/XI3/XI1/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM0 XROM/XI3/XI1/NET143 N_WL<26>_XROM/XI3/XI1/MM0_g
+ N_VSS_XROM/XI3/XI1/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM8 N_BL<0>_XROM/XI3/XI0/MM8_d N_WL<25>_XROM/XI3/XI0/MM8_g
+ N_VSS_XROM/XI3/XI0/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM0 XROM/XI3/XI0/NET143 N_WL<24>_XROM/XI3/XI0/MM0_g
+ N_VSS_XROM/XI3/XI0/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM8 N_BL<0>_XROM/XI2/XI3/MM8_d N_WL<23>_XROM/XI2/XI3/MM8_g
+ N_VSS_XROM/XI2/XI3/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM0 XROM/XI2/XI3/NET143 N_WL<22>_XROM/XI2/XI3/MM0_g
+ N_VSS_XROM/XI2/XI3/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM8 N_BL<0>_XROM/XI2/XI2/MM8_d N_WL<21>_XROM/XI2/XI2/MM8_g
+ N_VSS_XROM/XI2/XI2/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM0 XROM/XI2/XI2/NET143 N_WL<20>_XROM/XI2/XI2/MM0_g
+ N_VSS_XROM/XI2/XI2/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM8 N_BL<0>_XROM/XI2/XI1/MM8_d N_WL<19>_XROM/XI2/XI1/MM8_g
+ N_VSS_XROM/XI2/XI1/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM0 XROM/XI2/XI1/NET143 N_WL<18>_XROM/XI2/XI1/MM0_g
+ N_VSS_XROM/XI2/XI1/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM8 N_BL<0>_XROM/XI2/XI0/MM8_d N_WL<17>_XROM/XI2/XI0/MM8_g
+ N_VSS_XROM/XI2/XI0/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM0 XROM/XI2/XI0/NET143 N_WL<16>_XROM/XI2/XI0/MM0_g
+ N_VSS_XROM/XI2/XI0/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM9 XROM/XI3/XI3/NET107 N_WL<31>_XROM/XI3/XI3/MM9_g
+ N_VSS_XROM/XI3/XI3/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM1 N_BL<1>_XROM/XI3/XI3/MM1_d N_WL<30>_XROM/XI3/XI3/MM1_g
+ N_VSS_XROM/XI3/XI3/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM9 XROM/XI3/XI2/NET107 N_WL<29>_XROM/XI3/XI2/MM9_g
+ N_VSS_XROM/XI3/XI2/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM1 N_BL<1>_XROM/XI3/XI2/MM1_d N_WL<28>_XROM/XI3/XI2/MM1_g
+ N_VSS_XROM/XI3/XI2/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM9 XROM/XI3/XI1/NET107 N_WL<27>_XROM/XI3/XI1/MM9_g
+ N_VSS_XROM/XI3/XI1/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM1 N_BL<1>_XROM/XI3/XI1/MM1_d N_WL<26>_XROM/XI3/XI1/MM1_g
+ N_VSS_XROM/XI3/XI1/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM9 XROM/XI3/XI0/NET107 N_WL<25>_XROM/XI3/XI0/MM9_g
+ N_VSS_XROM/XI3/XI0/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM1 N_BL<1>_XROM/XI3/XI0/MM1_d N_WL<24>_XROM/XI3/XI0/MM1_g
+ N_VSS_XROM/XI3/XI0/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM9 XROM/XI2/XI3/NET107 N_WL<23>_XROM/XI2/XI3/MM9_g
+ N_VSS_XROM/XI2/XI3/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM1 N_BL<1>_XROM/XI2/XI3/MM1_d N_WL<22>_XROM/XI2/XI3/MM1_g
+ N_VSS_XROM/XI2/XI3/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM9 XROM/XI2/XI2/NET107 N_WL<21>_XROM/XI2/XI2/MM9_g
+ N_VSS_XROM/XI2/XI2/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM1 N_BL<1>_XROM/XI2/XI2/MM1_d N_WL<20>_XROM/XI2/XI2/MM1_g
+ N_VSS_XROM/XI2/XI2/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM9 XROM/XI2/XI1/NET107 N_WL<19>_XROM/XI2/XI1/MM9_g
+ N_VSS_XROM/XI2/XI1/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM1 N_BL<1>_XROM/XI2/XI1/MM1_d N_WL<18>_XROM/XI2/XI1/MM1_g
+ N_VSS_XROM/XI2/XI1/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM9 XROM/XI2/XI0/NET107 N_WL<17>_XROM/XI2/XI0/MM9_g
+ N_VSS_XROM/XI2/XI0/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM1 N_BL<1>_XROM/XI2/XI0/MM1_d N_WL<16>_XROM/XI2/XI0/MM1_g
+ N_VSS_XROM/XI2/XI0/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM10 N_BL<2>_XROM/XI3/XI3/MM10_d N_WL<31>_XROM/XI3/XI3/MM10_g
+ N_VSS_XROM/XI3/XI3/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM2 XROM/XI3/XI3/NET135 N_WL<30>_XROM/XI3/XI3/MM2_g
+ N_VSS_XROM/XI3/XI3/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM10 N_BL<2>_XROM/XI3/XI2/MM10_d N_WL<29>_XROM/XI3/XI2/MM10_g
+ N_VSS_XROM/XI3/XI2/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM2 XROM/XI3/XI2/NET135 N_WL<28>_XROM/XI3/XI2/MM2_g
+ N_VSS_XROM/XI3/XI2/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM10 N_BL<2>_XROM/XI3/XI1/MM10_d N_WL<27>_XROM/XI3/XI1/MM10_g
+ N_VSS_XROM/XI3/XI1/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM2 XROM/XI3/XI1/NET135 N_WL<26>_XROM/XI3/XI1/MM2_g
+ N_VSS_XROM/XI3/XI1/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM10 N_BL<2>_XROM/XI3/XI0/MM10_d N_WL<25>_XROM/XI3/XI0/MM10_g
+ N_VSS_XROM/XI3/XI0/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM2 XROM/XI3/XI0/NET135 N_WL<24>_XROM/XI3/XI0/MM2_g
+ N_VSS_XROM/XI3/XI0/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM10 N_BL<2>_XROM/XI2/XI3/MM10_d N_WL<23>_XROM/XI2/XI3/MM10_g
+ N_VSS_XROM/XI2/XI3/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM2 XROM/XI2/XI3/NET135 N_WL<22>_XROM/XI2/XI3/MM2_g
+ N_VSS_XROM/XI2/XI3/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM10 N_BL<2>_XROM/XI2/XI2/MM10_d N_WL<21>_XROM/XI2/XI2/MM10_g
+ N_VSS_XROM/XI2/XI2/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM2 XROM/XI2/XI2/NET135 N_WL<20>_XROM/XI2/XI2/MM2_g
+ N_VSS_XROM/XI2/XI2/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM10 N_BL<2>_XROM/XI2/XI1/MM10_d N_WL<19>_XROM/XI2/XI1/MM10_g
+ N_VSS_XROM/XI2/XI1/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM2 XROM/XI2/XI1/NET135 N_WL<18>_XROM/XI2/XI1/MM2_g
+ N_VSS_XROM/XI2/XI1/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM10 N_BL<2>_XROM/XI2/XI0/MM10_d N_WL<17>_XROM/XI2/XI0/MM10_g
+ N_VSS_XROM/XI2/XI0/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM2 XROM/XI2/XI0/NET135 N_WL<16>_XROM/XI2/XI0/MM2_g
+ N_VSS_XROM/XI2/XI0/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM11 XROM/XI3/XI3/NET99 N_WL<31>_XROM/XI3/XI3/MM11_g
+ N_VSS_XROM/XI3/XI3/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM3 N_BL<3>_XROM/XI3/XI3/MM3_d N_WL<30>_XROM/XI3/XI3/MM3_g
+ N_VSS_XROM/XI3/XI3/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM11 XROM/XI3/XI2/NET99 N_WL<29>_XROM/XI3/XI2/MM11_g
+ N_VSS_XROM/XI3/XI2/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM3 N_BL<3>_XROM/XI3/XI2/MM3_d N_WL<28>_XROM/XI3/XI2/MM3_g
+ N_VSS_XROM/XI3/XI2/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM11 XROM/XI3/XI1/NET99 N_WL<27>_XROM/XI3/XI1/MM11_g
+ N_VSS_XROM/XI3/XI1/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM3 N_BL<3>_XROM/XI3/XI1/MM3_d N_WL<26>_XROM/XI3/XI1/MM3_g
+ N_VSS_XROM/XI3/XI1/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM11 XROM/XI3/XI0/NET99 N_WL<25>_XROM/XI3/XI0/MM11_g
+ N_VSS_XROM/XI3/XI0/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM3 N_BL<3>_XROM/XI3/XI0/MM3_d N_WL<24>_XROM/XI3/XI0/MM3_g
+ N_VSS_XROM/XI3/XI0/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM11 XROM/XI2/XI3/NET99 N_WL<23>_XROM/XI2/XI3/MM11_g
+ N_VSS_XROM/XI2/XI3/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM3 N_BL<3>_XROM/XI2/XI3/MM3_d N_WL<22>_XROM/XI2/XI3/MM3_g
+ N_VSS_XROM/XI2/XI3/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM11 XROM/XI2/XI2/NET99 N_WL<21>_XROM/XI2/XI2/MM11_g
+ N_VSS_XROM/XI2/XI2/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM3 N_BL<3>_XROM/XI2/XI2/MM3_d N_WL<20>_XROM/XI2/XI2/MM3_g
+ N_VSS_XROM/XI2/XI2/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM11 XROM/XI2/XI1/NET99 N_WL<19>_XROM/XI2/XI1/MM11_g
+ N_VSS_XROM/XI2/XI1/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM3 N_BL<3>_XROM/XI2/XI1/MM3_d N_WL<18>_XROM/XI2/XI1/MM3_g
+ N_VSS_XROM/XI2/XI1/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM11 XROM/XI2/XI0/NET99 N_WL<17>_XROM/XI2/XI0/MM11_g
+ N_VSS_XROM/XI2/XI0/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM3 N_BL<3>_XROM/XI2/XI0/MM3_d N_WL<16>_XROM/XI2/XI0/MM3_g
+ N_VSS_XROM/XI2/XI0/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM12 N_BL<4>_XROM/XI3/XI3/MM12_d N_WL<31>_XROM/XI3/XI3/MM12_g
+ N_VSS_XROM/XI3/XI3/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM4 XROM/XI3/XI3/NET127 N_WL<30>_XROM/XI3/XI3/MM4_g
+ N_VSS_XROM/XI3/XI3/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM12 N_BL<4>_XROM/XI3/XI2/MM12_d N_WL<29>_XROM/XI3/XI2/MM12_g
+ N_VSS_XROM/XI3/XI2/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM4 XROM/XI3/XI2/NET127 N_WL<28>_XROM/XI3/XI2/MM4_g
+ N_VSS_XROM/XI3/XI2/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM12 N_BL<4>_XROM/XI3/XI1/MM12_d N_WL<27>_XROM/XI3/XI1/MM12_g
+ N_VSS_XROM/XI3/XI1/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM4 XROM/XI3/XI1/NET127 N_WL<26>_XROM/XI3/XI1/MM4_g
+ N_VSS_XROM/XI3/XI1/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM12 N_BL<4>_XROM/XI3/XI0/MM12_d N_WL<25>_XROM/XI3/XI0/MM12_g
+ N_VSS_XROM/XI3/XI0/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM4 XROM/XI3/XI0/NET127 N_WL<24>_XROM/XI3/XI0/MM4_g
+ N_VSS_XROM/XI3/XI0/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM12 N_BL<4>_XROM/XI2/XI3/MM12_d N_WL<23>_XROM/XI2/XI3/MM12_g
+ N_VSS_XROM/XI2/XI3/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM4 XROM/XI2/XI3/NET127 N_WL<22>_XROM/XI2/XI3/MM4_g
+ N_VSS_XROM/XI2/XI3/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM12 N_BL<4>_XROM/XI2/XI2/MM12_d N_WL<21>_XROM/XI2/XI2/MM12_g
+ N_VSS_XROM/XI2/XI2/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM4 XROM/XI2/XI2/NET127 N_WL<20>_XROM/XI2/XI2/MM4_g
+ N_VSS_XROM/XI2/XI2/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM12 N_BL<4>_XROM/XI2/XI1/MM12_d N_WL<19>_XROM/XI2/XI1/MM12_g
+ N_VSS_XROM/XI2/XI1/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM4 XROM/XI2/XI1/NET127 N_WL<18>_XROM/XI2/XI1/MM4_g
+ N_VSS_XROM/XI2/XI1/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM12 N_BL<4>_XROM/XI2/XI0/MM12_d N_WL<17>_XROM/XI2/XI0/MM12_g
+ N_VSS_XROM/XI2/XI0/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM4 XROM/XI2/XI0/NET127 N_WL<16>_XROM/XI2/XI0/MM4_g
+ N_VSS_XROM/XI2/XI0/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM13 XROM/XI3/XI3/NET91 N_WL<31>_XROM/XI3/XI3/MM13_g
+ N_VSS_XROM/XI3/XI3/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM5 N_BL<5>_XROM/XI3/XI3/MM5_d N_WL<30>_XROM/XI3/XI3/MM5_g
+ N_VSS_XROM/XI3/XI3/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM13 XROM/XI3/XI2/NET91 N_WL<29>_XROM/XI3/XI2/MM13_g
+ N_VSS_XROM/XI3/XI2/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM5 N_BL<5>_XROM/XI3/XI2/MM5_d N_WL<28>_XROM/XI3/XI2/MM5_g
+ N_VSS_XROM/XI3/XI2/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM13 XROM/XI3/XI1/NET91 N_WL<27>_XROM/XI3/XI1/MM13_g
+ N_VSS_XROM/XI3/XI1/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM5 N_BL<5>_XROM/XI3/XI1/MM5_d N_WL<26>_XROM/XI3/XI1/MM5_g
+ N_VSS_XROM/XI3/XI1/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM13 XROM/XI3/XI0/NET91 N_WL<25>_XROM/XI3/XI0/MM13_g
+ N_VSS_XROM/XI3/XI0/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM5 N_BL<5>_XROM/XI3/XI0/MM5_d N_WL<24>_XROM/XI3/XI0/MM5_g
+ N_VSS_XROM/XI3/XI0/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM13 XROM/XI2/XI3/NET91 N_WL<23>_XROM/XI2/XI3/MM13_g
+ N_VSS_XROM/XI2/XI3/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM5 N_BL<5>_XROM/XI2/XI3/MM5_d N_WL<22>_XROM/XI2/XI3/MM5_g
+ N_VSS_XROM/XI2/XI3/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM13 XROM/XI2/XI2/NET91 N_WL<21>_XROM/XI2/XI2/MM13_g
+ N_VSS_XROM/XI2/XI2/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM5 N_BL<5>_XROM/XI2/XI2/MM5_d N_WL<20>_XROM/XI2/XI2/MM5_g
+ N_VSS_XROM/XI2/XI2/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM13 XROM/XI2/XI1/NET91 N_WL<19>_XROM/XI2/XI1/MM13_g
+ N_VSS_XROM/XI2/XI1/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM5 N_BL<5>_XROM/XI2/XI1/MM5_d N_WL<18>_XROM/XI2/XI1/MM5_g
+ N_VSS_XROM/XI2/XI1/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM13 XROM/XI2/XI0/NET91 N_WL<17>_XROM/XI2/XI0/MM13_g
+ N_VSS_XROM/XI2/XI0/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM5 N_BL<5>_XROM/XI2/XI0/MM5_d N_WL<16>_XROM/XI2/XI0/MM5_g
+ N_VSS_XROM/XI2/XI0/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM14 N_BL<6>_XROM/XI3/XI3/MM14_d N_WL<31>_XROM/XI3/XI3/MM14_g
+ N_VSS_XROM/XI3/XI3/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM6 XROM/XI3/XI3/NET119 N_WL<30>_XROM/XI3/XI3/MM6_g
+ N_VSS_XROM/XI3/XI3/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM14 N_BL<6>_XROM/XI3/XI2/MM14_d N_WL<29>_XROM/XI3/XI2/MM14_g
+ N_VSS_XROM/XI3/XI2/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM6 XROM/XI3/XI2/NET119 N_WL<28>_XROM/XI3/XI2/MM6_g
+ N_VSS_XROM/XI3/XI2/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM14 N_BL<6>_XROM/XI3/XI1/MM14_d N_WL<27>_XROM/XI3/XI1/MM14_g
+ N_VSS_XROM/XI3/XI1/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM6 XROM/XI3/XI1/NET119 N_WL<26>_XROM/XI3/XI1/MM6_g
+ N_VSS_XROM/XI3/XI1/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM14 N_BL<6>_XROM/XI3/XI0/MM14_d N_WL<25>_XROM/XI3/XI0/MM14_g
+ N_VSS_XROM/XI3/XI0/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM6 XROM/XI3/XI0/NET119 N_WL<24>_XROM/XI3/XI0/MM6_g
+ N_VSS_XROM/XI3/XI0/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM14 N_BL<6>_XROM/XI2/XI3/MM14_d N_WL<23>_XROM/XI2/XI3/MM14_g
+ N_VSS_XROM/XI2/XI3/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM6 XROM/XI2/XI3/NET119 N_WL<22>_XROM/XI2/XI3/MM6_g
+ N_VSS_XROM/XI2/XI3/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM14 N_BL<6>_XROM/XI2/XI2/MM14_d N_WL<21>_XROM/XI2/XI2/MM14_g
+ N_VSS_XROM/XI2/XI2/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM6 XROM/XI2/XI2/NET119 N_WL<20>_XROM/XI2/XI2/MM6_g
+ N_VSS_XROM/XI2/XI2/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM14 N_BL<6>_XROM/XI2/XI1/MM14_d N_WL<19>_XROM/XI2/XI1/MM14_g
+ N_VSS_XROM/XI2/XI1/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM6 XROM/XI2/XI1/NET119 N_WL<18>_XROM/XI2/XI1/MM6_g
+ N_VSS_XROM/XI2/XI1/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM14 N_BL<6>_XROM/XI2/XI0/MM14_d N_WL<17>_XROM/XI2/XI0/MM14_g
+ N_VSS_XROM/XI2/XI0/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM6 XROM/XI2/XI0/NET119 N_WL<16>_XROM/XI2/XI0/MM6_g
+ N_VSS_XROM/XI2/XI0/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM15 XROM/XI3/XI3/NET83 N_WL<31>_XROM/XI3/XI3/MM15_g
+ N_VSS_XROM/XI3/XI3/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI3/MM7 N_BL<7>_XROM/XI3/XI3/MM7_d N_WL<30>_XROM/XI3/XI3/MM7_g
+ N_VSS_XROM/XI3/XI3/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM15 XROM/XI3/XI2/NET83 N_WL<29>_XROM/XI3/XI2/MM15_g
+ N_VSS_XROM/XI3/XI2/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI2/MM7 N_BL<7>_XROM/XI3/XI2/MM7_d N_WL<28>_XROM/XI3/XI2/MM7_g
+ N_VSS_XROM/XI3/XI2/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM15 XROM/XI3/XI1/NET83 N_WL<27>_XROM/XI3/XI1/MM15_g
+ N_VSS_XROM/XI3/XI1/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI1/MM7 N_BL<7>_XROM/XI3/XI1/MM7_d N_WL<26>_XROM/XI3/XI1/MM7_g
+ N_VSS_XROM/XI3/XI1/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM15 XROM/XI3/XI0/NET83 N_WL<25>_XROM/XI3/XI0/MM15_g
+ N_VSS_XROM/XI3/XI0/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI0/MM7 N_BL<7>_XROM/XI3/XI0/MM7_d N_WL<24>_XROM/XI3/XI0/MM7_g
+ N_VSS_XROM/XI3/XI0/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM15 XROM/XI2/XI3/NET83 N_WL<23>_XROM/XI2/XI3/MM15_g
+ N_VSS_XROM/XI2/XI3/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI3/MM7 N_BL<7>_XROM/XI2/XI3/MM7_d N_WL<22>_XROM/XI2/XI3/MM7_g
+ N_VSS_XROM/XI2/XI3/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM15 XROM/XI2/XI2/NET83 N_WL<21>_XROM/XI2/XI2/MM15_g
+ N_VSS_XROM/XI2/XI2/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI2/MM7 N_BL<7>_XROM/XI2/XI2/MM7_d N_WL<20>_XROM/XI2/XI2/MM7_g
+ N_VSS_XROM/XI2/XI2/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM15 XROM/XI2/XI1/NET83 N_WL<19>_XROM/XI2/XI1/MM15_g
+ N_VSS_XROM/XI2/XI1/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI1/MM7 N_BL<7>_XROM/XI2/XI1/MM7_d N_WL<18>_XROM/XI2/XI1/MM7_g
+ N_VSS_XROM/XI2/XI1/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM15 XROM/XI2/XI0/NET83 N_WL<17>_XROM/XI2/XI0/MM15_g
+ N_VSS_XROM/XI2/XI0/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI0/MM7 N_BL<7>_XROM/XI2/XI0/MM7_d N_WL<16>_XROM/XI2/XI0/MM7_g
+ N_VSS_XROM/XI2/XI0/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM8 N_BL<8>_XROM/XI3/XI7/MM8_d N_WL<31>_XROM/XI3/XI7/MM8_g
+ N_VSS_XROM/XI3/XI7/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM0 XROM/XI3/XI7/NET143 N_WL<30>_XROM/XI3/XI7/MM0_g
+ N_VSS_XROM/XI3/XI7/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM8 N_BL<8>_XROM/XI3/XI6/MM8_d N_WL<29>_XROM/XI3/XI6/MM8_g
+ N_VSS_XROM/XI3/XI6/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM0 XROM/XI3/XI6/NET143 N_WL<28>_XROM/XI3/XI6/MM0_g
+ N_VSS_XROM/XI3/XI6/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM8 N_BL<8>_XROM/XI3/XI5/MM8_d N_WL<27>_XROM/XI3/XI5/MM8_g
+ N_VSS_XROM/XI3/XI5/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM0 XROM/XI3/XI5/NET143 N_WL<26>_XROM/XI3/XI5/MM0_g
+ N_VSS_XROM/XI3/XI5/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM8 N_BL<8>_XROM/XI3/XI4/MM8_d N_WL<25>_XROM/XI3/XI4/MM8_g
+ N_VSS_XROM/XI3/XI4/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM0 XROM/XI3/XI4/NET143 N_WL<24>_XROM/XI3/XI4/MM0_g
+ N_VSS_XROM/XI3/XI4/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM8 N_BL<8>_XROM/XI2/XI7/MM8_d N_WL<23>_XROM/XI2/XI7/MM8_g
+ N_VSS_XROM/XI2/XI7/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM0 XROM/XI2/XI7/NET143 N_WL<22>_XROM/XI2/XI7/MM0_g
+ N_VSS_XROM/XI2/XI7/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM8 N_BL<8>_XROM/XI2/XI6/MM8_d N_WL<21>_XROM/XI2/XI6/MM8_g
+ N_VSS_XROM/XI2/XI6/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM0 XROM/XI2/XI6/NET143 N_WL<20>_XROM/XI2/XI6/MM0_g
+ N_VSS_XROM/XI2/XI6/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM8 N_BL<8>_XROM/XI2/XI5/MM8_d N_WL<19>_XROM/XI2/XI5/MM8_g
+ N_VSS_XROM/XI2/XI5/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM0 XROM/XI2/XI5/NET143 N_WL<18>_XROM/XI2/XI5/MM0_g
+ N_VSS_XROM/XI2/XI5/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM8 N_BL<8>_XROM/XI2/XI4/MM8_d N_WL<17>_XROM/XI2/XI4/MM8_g
+ N_VSS_XROM/XI2/XI4/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM0 XROM/XI2/XI4/NET143 N_WL<16>_XROM/XI2/XI4/MM0_g
+ N_VSS_XROM/XI2/XI4/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM9 XROM/XI3/XI7/NET107 N_WL<31>_XROM/XI3/XI7/MM9_g
+ N_VSS_XROM/XI3/XI7/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM1 N_BL<9>_XROM/XI3/XI7/MM1_d N_WL<30>_XROM/XI3/XI7/MM1_g
+ N_VSS_XROM/XI3/XI7/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM9 XROM/XI3/XI6/NET107 N_WL<29>_XROM/XI3/XI6/MM9_g
+ N_VSS_XROM/XI3/XI6/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM1 N_BL<9>_XROM/XI3/XI6/MM1_d N_WL<28>_XROM/XI3/XI6/MM1_g
+ N_VSS_XROM/XI3/XI6/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM9 XROM/XI3/XI5/NET107 N_WL<27>_XROM/XI3/XI5/MM9_g
+ N_VSS_XROM/XI3/XI5/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM1 N_BL<9>_XROM/XI3/XI5/MM1_d N_WL<26>_XROM/XI3/XI5/MM1_g
+ N_VSS_XROM/XI3/XI5/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM9 XROM/XI3/XI4/NET107 N_WL<25>_XROM/XI3/XI4/MM9_g
+ N_VSS_XROM/XI3/XI4/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM1 N_BL<9>_XROM/XI3/XI4/MM1_d N_WL<24>_XROM/XI3/XI4/MM1_g
+ N_VSS_XROM/XI3/XI4/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM9 XROM/XI2/XI7/NET107 N_WL<23>_XROM/XI2/XI7/MM9_g
+ N_VSS_XROM/XI2/XI7/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM1 N_BL<9>_XROM/XI2/XI7/MM1_d N_WL<22>_XROM/XI2/XI7/MM1_g
+ N_VSS_XROM/XI2/XI7/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM9 XROM/XI2/XI6/NET107 N_WL<21>_XROM/XI2/XI6/MM9_g
+ N_VSS_XROM/XI2/XI6/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM1 N_BL<9>_XROM/XI2/XI6/MM1_d N_WL<20>_XROM/XI2/XI6/MM1_g
+ N_VSS_XROM/XI2/XI6/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM9 XROM/XI2/XI5/NET107 N_WL<19>_XROM/XI2/XI5/MM9_g
+ N_VSS_XROM/XI2/XI5/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM1 N_BL<9>_XROM/XI2/XI5/MM1_d N_WL<18>_XROM/XI2/XI5/MM1_g
+ N_VSS_XROM/XI2/XI5/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM9 XROM/XI2/XI4/NET107 N_WL<17>_XROM/XI2/XI4/MM9_g
+ N_VSS_XROM/XI2/XI4/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM1 N_BL<9>_XROM/XI2/XI4/MM1_d N_WL<16>_XROM/XI2/XI4/MM1_g
+ N_VSS_XROM/XI2/XI4/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM10 N_BL<10>_XROM/XI3/XI7/MM10_d N_WL<31>_XROM/XI3/XI7/MM10_g
+ N_VSS_XROM/XI3/XI7/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM2 XROM/XI3/XI7/NET135 N_WL<30>_XROM/XI3/XI7/MM2_g
+ N_VSS_XROM/XI3/XI7/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM10 N_BL<10>_XROM/XI3/XI6/MM10_d N_WL<29>_XROM/XI3/XI6/MM10_g
+ N_VSS_XROM/XI3/XI6/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM2 XROM/XI3/XI6/NET135 N_WL<28>_XROM/XI3/XI6/MM2_g
+ N_VSS_XROM/XI3/XI6/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM10 N_BL<10>_XROM/XI3/XI5/MM10_d N_WL<27>_XROM/XI3/XI5/MM10_g
+ N_VSS_XROM/XI3/XI5/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM2 XROM/XI3/XI5/NET135 N_WL<26>_XROM/XI3/XI5/MM2_g
+ N_VSS_XROM/XI3/XI5/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM10 N_BL<10>_XROM/XI3/XI4/MM10_d N_WL<25>_XROM/XI3/XI4/MM10_g
+ N_VSS_XROM/XI3/XI4/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM2 XROM/XI3/XI4/NET135 N_WL<24>_XROM/XI3/XI4/MM2_g
+ N_VSS_XROM/XI3/XI4/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM10 N_BL<10>_XROM/XI2/XI7/MM10_d N_WL<23>_XROM/XI2/XI7/MM10_g
+ N_VSS_XROM/XI2/XI7/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM2 XROM/XI2/XI7/NET135 N_WL<22>_XROM/XI2/XI7/MM2_g
+ N_VSS_XROM/XI2/XI7/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM10 N_BL<10>_XROM/XI2/XI6/MM10_d N_WL<21>_XROM/XI2/XI6/MM10_g
+ N_VSS_XROM/XI2/XI6/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM2 XROM/XI2/XI6/NET135 N_WL<20>_XROM/XI2/XI6/MM2_g
+ N_VSS_XROM/XI2/XI6/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM10 N_BL<10>_XROM/XI2/XI5/MM10_d N_WL<19>_XROM/XI2/XI5/MM10_g
+ N_VSS_XROM/XI2/XI5/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM2 XROM/XI2/XI5/NET135 N_WL<18>_XROM/XI2/XI5/MM2_g
+ N_VSS_XROM/XI2/XI5/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM10 N_BL<10>_XROM/XI2/XI4/MM10_d N_WL<17>_XROM/XI2/XI4/MM10_g
+ N_VSS_XROM/XI2/XI4/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM2 XROM/XI2/XI4/NET135 N_WL<16>_XROM/XI2/XI4/MM2_g
+ N_VSS_XROM/XI2/XI4/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM11 XROM/XI3/XI7/NET99 N_WL<31>_XROM/XI3/XI7/MM11_g
+ N_VSS_XROM/XI3/XI7/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM3 N_BL<11>_XROM/XI3/XI7/MM3_d N_WL<30>_XROM/XI3/XI7/MM3_g
+ N_VSS_XROM/XI3/XI7/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM11 XROM/XI3/XI6/NET99 N_WL<29>_XROM/XI3/XI6/MM11_g
+ N_VSS_XROM/XI3/XI6/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM3 N_BL<11>_XROM/XI3/XI6/MM3_d N_WL<28>_XROM/XI3/XI6/MM3_g
+ N_VSS_XROM/XI3/XI6/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM11 XROM/XI3/XI5/NET99 N_WL<27>_XROM/XI3/XI5/MM11_g
+ N_VSS_XROM/XI3/XI5/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM3 N_BL<11>_XROM/XI3/XI5/MM3_d N_WL<26>_XROM/XI3/XI5/MM3_g
+ N_VSS_XROM/XI3/XI5/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM11 XROM/XI3/XI4/NET99 N_WL<25>_XROM/XI3/XI4/MM11_g
+ N_VSS_XROM/XI3/XI4/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM3 N_BL<11>_XROM/XI3/XI4/MM3_d N_WL<24>_XROM/XI3/XI4/MM3_g
+ N_VSS_XROM/XI3/XI4/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM11 XROM/XI2/XI7/NET99 N_WL<23>_XROM/XI2/XI7/MM11_g
+ N_VSS_XROM/XI2/XI7/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM3 N_BL<11>_XROM/XI2/XI7/MM3_d N_WL<22>_XROM/XI2/XI7/MM3_g
+ N_VSS_XROM/XI2/XI7/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM11 XROM/XI2/XI6/NET99 N_WL<21>_XROM/XI2/XI6/MM11_g
+ N_VSS_XROM/XI2/XI6/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM3 N_BL<11>_XROM/XI2/XI6/MM3_d N_WL<20>_XROM/XI2/XI6/MM3_g
+ N_VSS_XROM/XI2/XI6/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM11 XROM/XI2/XI5/NET99 N_WL<19>_XROM/XI2/XI5/MM11_g
+ N_VSS_XROM/XI2/XI5/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM3 N_BL<11>_XROM/XI2/XI5/MM3_d N_WL<18>_XROM/XI2/XI5/MM3_g
+ N_VSS_XROM/XI2/XI5/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM11 XROM/XI2/XI4/NET99 N_WL<17>_XROM/XI2/XI4/MM11_g
+ N_VSS_XROM/XI2/XI4/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM3 N_BL<11>_XROM/XI2/XI4/MM3_d N_WL<16>_XROM/XI2/XI4/MM3_g
+ N_VSS_XROM/XI2/XI4/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM12 N_BL<12>_XROM/XI3/XI7/MM12_d N_WL<31>_XROM/XI3/XI7/MM12_g
+ N_VSS_XROM/XI3/XI7/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM4 XROM/XI3/XI7/NET127 N_WL<30>_XROM/XI3/XI7/MM4_g
+ N_VSS_XROM/XI3/XI7/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM12 N_BL<12>_XROM/XI3/XI6/MM12_d N_WL<29>_XROM/XI3/XI6/MM12_g
+ N_VSS_XROM/XI3/XI6/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM4 XROM/XI3/XI6/NET127 N_WL<28>_XROM/XI3/XI6/MM4_g
+ N_VSS_XROM/XI3/XI6/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM12 N_BL<12>_XROM/XI3/XI5/MM12_d N_WL<27>_XROM/XI3/XI5/MM12_g
+ N_VSS_XROM/XI3/XI5/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM4 XROM/XI3/XI5/NET127 N_WL<26>_XROM/XI3/XI5/MM4_g
+ N_VSS_XROM/XI3/XI5/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM12 N_BL<12>_XROM/XI3/XI4/MM12_d N_WL<25>_XROM/XI3/XI4/MM12_g
+ N_VSS_XROM/XI3/XI4/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM4 XROM/XI3/XI4/NET127 N_WL<24>_XROM/XI3/XI4/MM4_g
+ N_VSS_XROM/XI3/XI4/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM12 N_BL<12>_XROM/XI2/XI7/MM12_d N_WL<23>_XROM/XI2/XI7/MM12_g
+ N_VSS_XROM/XI2/XI7/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM4 XROM/XI2/XI7/NET127 N_WL<22>_XROM/XI2/XI7/MM4_g
+ N_VSS_XROM/XI2/XI7/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM12 N_BL<12>_XROM/XI2/XI6/MM12_d N_WL<21>_XROM/XI2/XI6/MM12_g
+ N_VSS_XROM/XI2/XI6/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM4 XROM/XI2/XI6/NET127 N_WL<20>_XROM/XI2/XI6/MM4_g
+ N_VSS_XROM/XI2/XI6/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM12 N_BL<12>_XROM/XI2/XI5/MM12_d N_WL<19>_XROM/XI2/XI5/MM12_g
+ N_VSS_XROM/XI2/XI5/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM4 XROM/XI2/XI5/NET127 N_WL<18>_XROM/XI2/XI5/MM4_g
+ N_VSS_XROM/XI2/XI5/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM12 N_BL<12>_XROM/XI2/XI4/MM12_d N_WL<17>_XROM/XI2/XI4/MM12_g
+ N_VSS_XROM/XI2/XI4/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM4 XROM/XI2/XI4/NET127 N_WL<16>_XROM/XI2/XI4/MM4_g
+ N_VSS_XROM/XI2/XI4/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM13 XROM/XI3/XI7/NET91 N_WL<31>_XROM/XI3/XI7/MM13_g
+ N_VSS_XROM/XI3/XI7/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM5 N_BL<13>_XROM/XI3/XI7/MM5_d N_WL<30>_XROM/XI3/XI7/MM5_g
+ N_VSS_XROM/XI3/XI7/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM13 XROM/XI3/XI6/NET91 N_WL<29>_XROM/XI3/XI6/MM13_g
+ N_VSS_XROM/XI3/XI6/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM5 N_BL<13>_XROM/XI3/XI6/MM5_d N_WL<28>_XROM/XI3/XI6/MM5_g
+ N_VSS_XROM/XI3/XI6/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM13 XROM/XI3/XI5/NET91 N_WL<27>_XROM/XI3/XI5/MM13_g
+ N_VSS_XROM/XI3/XI5/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM5 N_BL<13>_XROM/XI3/XI5/MM5_d N_WL<26>_XROM/XI3/XI5/MM5_g
+ N_VSS_XROM/XI3/XI5/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM13 XROM/XI3/XI4/NET91 N_WL<25>_XROM/XI3/XI4/MM13_g
+ N_VSS_XROM/XI3/XI4/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM5 N_BL<13>_XROM/XI3/XI4/MM5_d N_WL<24>_XROM/XI3/XI4/MM5_g
+ N_VSS_XROM/XI3/XI4/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM13 XROM/XI2/XI7/NET91 N_WL<23>_XROM/XI2/XI7/MM13_g
+ N_VSS_XROM/XI2/XI7/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM5 N_BL<13>_XROM/XI2/XI7/MM5_d N_WL<22>_XROM/XI2/XI7/MM5_g
+ N_VSS_XROM/XI2/XI7/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM13 XROM/XI2/XI6/NET91 N_WL<21>_XROM/XI2/XI6/MM13_g
+ N_VSS_XROM/XI2/XI6/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM5 N_BL<13>_XROM/XI2/XI6/MM5_d N_WL<20>_XROM/XI2/XI6/MM5_g
+ N_VSS_XROM/XI2/XI6/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM13 XROM/XI2/XI5/NET91 N_WL<19>_XROM/XI2/XI5/MM13_g
+ N_VSS_XROM/XI2/XI5/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM5 N_BL<13>_XROM/XI2/XI5/MM5_d N_WL<18>_XROM/XI2/XI5/MM5_g
+ N_VSS_XROM/XI2/XI5/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM13 XROM/XI2/XI4/NET91 N_WL<17>_XROM/XI2/XI4/MM13_g
+ N_VSS_XROM/XI2/XI4/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM5 N_BL<13>_XROM/XI2/XI4/MM5_d N_WL<16>_XROM/XI2/XI4/MM5_g
+ N_VSS_XROM/XI2/XI4/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM14 N_BL<14>_XROM/XI3/XI7/MM14_d N_WL<31>_XROM/XI3/XI7/MM14_g
+ N_VSS_XROM/XI3/XI7/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM6 XROM/XI3/XI7/NET119 N_WL<30>_XROM/XI3/XI7/MM6_g
+ N_VSS_XROM/XI3/XI7/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM14 N_BL<14>_XROM/XI3/XI6/MM14_d N_WL<29>_XROM/XI3/XI6/MM14_g
+ N_VSS_XROM/XI3/XI6/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM6 XROM/XI3/XI6/NET119 N_WL<28>_XROM/XI3/XI6/MM6_g
+ N_VSS_XROM/XI3/XI6/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM14 N_BL<14>_XROM/XI3/XI5/MM14_d N_WL<27>_XROM/XI3/XI5/MM14_g
+ N_VSS_XROM/XI3/XI5/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM6 XROM/XI3/XI5/NET119 N_WL<26>_XROM/XI3/XI5/MM6_g
+ N_VSS_XROM/XI3/XI5/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM14 N_BL<14>_XROM/XI3/XI4/MM14_d N_WL<25>_XROM/XI3/XI4/MM14_g
+ N_VSS_XROM/XI3/XI4/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM6 XROM/XI3/XI4/NET119 N_WL<24>_XROM/XI3/XI4/MM6_g
+ N_VSS_XROM/XI3/XI4/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM14 N_BL<14>_XROM/XI2/XI7/MM14_d N_WL<23>_XROM/XI2/XI7/MM14_g
+ N_VSS_XROM/XI2/XI7/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM6 XROM/XI2/XI7/NET119 N_WL<22>_XROM/XI2/XI7/MM6_g
+ N_VSS_XROM/XI2/XI7/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM14 N_BL<14>_XROM/XI2/XI6/MM14_d N_WL<21>_XROM/XI2/XI6/MM14_g
+ N_VSS_XROM/XI2/XI6/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM6 XROM/XI2/XI6/NET119 N_WL<20>_XROM/XI2/XI6/MM6_g
+ N_VSS_XROM/XI2/XI6/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM14 N_BL<14>_XROM/XI2/XI5/MM14_d N_WL<19>_XROM/XI2/XI5/MM14_g
+ N_VSS_XROM/XI2/XI5/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM6 XROM/XI2/XI5/NET119 N_WL<18>_XROM/XI2/XI5/MM6_g
+ N_VSS_XROM/XI2/XI5/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM14 N_BL<14>_XROM/XI2/XI4/MM14_d N_WL<17>_XROM/XI2/XI4/MM14_g
+ N_VSS_XROM/XI2/XI4/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM6 XROM/XI2/XI4/NET119 N_WL<16>_XROM/XI2/XI4/MM6_g
+ N_VSS_XROM/XI2/XI4/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM15 XROM/XI3/XI7/NET83 N_WL<31>_XROM/XI3/XI7/MM15_g
+ N_VSS_XROM/XI3/XI7/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI7/MM7 N_BL<15>_XROM/XI3/XI7/MM7_d N_WL<30>_XROM/XI3/XI7/MM7_g
+ N_VSS_XROM/XI3/XI7/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM15 XROM/XI3/XI6/NET83 N_WL<29>_XROM/XI3/XI6/MM15_g
+ N_VSS_XROM/XI3/XI6/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI6/MM7 N_BL<15>_XROM/XI3/XI6/MM7_d N_WL<28>_XROM/XI3/XI6/MM7_g
+ N_VSS_XROM/XI3/XI6/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM15 XROM/XI3/XI5/NET83 N_WL<27>_XROM/XI3/XI5/MM15_g
+ N_VSS_XROM/XI3/XI5/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI5/MM7 N_BL<15>_XROM/XI3/XI5/MM7_d N_WL<26>_XROM/XI3/XI5/MM7_g
+ N_VSS_XROM/XI3/XI5/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM15 XROM/XI3/XI4/NET83 N_WL<25>_XROM/XI3/XI4/MM15_g
+ N_VSS_XROM/XI3/XI4/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI3/XI4/MM7 N_BL<15>_XROM/XI3/XI4/MM7_d N_WL<24>_XROM/XI3/XI4/MM7_g
+ N_VSS_XROM/XI3/XI4/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM15 XROM/XI2/XI7/NET83 N_WL<23>_XROM/XI2/XI7/MM15_g
+ N_VSS_XROM/XI2/XI7/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI7/MM7 N_BL<15>_XROM/XI2/XI7/MM7_d N_WL<22>_XROM/XI2/XI7/MM7_g
+ N_VSS_XROM/XI2/XI7/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM15 XROM/XI2/XI6/NET83 N_WL<21>_XROM/XI2/XI6/MM15_g
+ N_VSS_XROM/XI2/XI6/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI6/MM7 N_BL<15>_XROM/XI2/XI6/MM7_d N_WL<20>_XROM/XI2/XI6/MM7_g
+ N_VSS_XROM/XI2/XI6/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM15 XROM/XI2/XI5/NET83 N_WL<19>_XROM/XI2/XI5/MM15_g
+ N_VSS_XROM/XI2/XI5/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI5/MM7 N_BL<15>_XROM/XI2/XI5/MM7_d N_WL<18>_XROM/XI2/XI5/MM7_g
+ N_VSS_XROM/XI2/XI5/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM15 XROM/XI2/XI4/NET83 N_WL<17>_XROM/XI2/XI4/MM15_g
+ N_VSS_XROM/XI2/XI4/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI2/XI4/MM7 N_BL<15>_XROM/XI2/XI4/MM7_d N_WL<16>_XROM/XI2/XI4/MM7_g
+ N_VSS_XROM/XI2/XI4/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM8 N_BL<0>_XROM/XI1/XI3/MM8_d N_WL<15>_XROM/XI1/XI3/MM8_g
+ N_VSS_XROM/XI1/XI3/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM0 XROM/XI1/XI3/NET143 N_WL<14>_XROM/XI1/XI3/MM0_g
+ N_VSS_XROM/XI1/XI3/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM8 N_BL<0>_XROM/XI1/XI2/MM8_d N_WL<13>_XROM/XI1/XI2/MM8_g
+ N_VSS_XROM/XI1/XI2/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM0 XROM/XI1/XI2/NET143 N_WL<12>_XROM/XI1/XI2/MM0_g
+ N_VSS_XROM/XI1/XI2/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM8 N_BL<0>_XROM/XI1/XI1/MM8_d N_WL<11>_XROM/XI1/XI1/MM8_g
+ N_VSS_XROM/XI1/XI1/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM0 XROM/XI1/XI1/NET143 N_WL<10>_XROM/XI1/XI1/MM0_g
+ N_VSS_XROM/XI1/XI1/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM8 N_BL<0>_XROM/XI1/XI0/MM8_d N_WL<9>_XROM/XI1/XI0/MM8_g
+ N_VSS_XROM/XI1/XI0/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM0 XROM/XI1/XI0/NET143 N_WL<8>_XROM/XI1/XI0/MM0_g
+ N_VSS_XROM/XI1/XI0/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM8 N_BL<0>_XROM/XI0/XI3/MM8_d N_WL<7>_XROM/XI0/XI3/MM8_g
+ N_VSS_XROM/XI0/XI3/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM0 XROM/XI0/XI3/NET143 N_WL<6>_XROM/XI0/XI3/MM0_g
+ N_VSS_XROM/XI0/XI3/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM8 N_BL<0>_XROM/XI0/XI2/MM8_d N_WL<5>_XROM/XI0/XI2/MM8_g
+ N_VSS_XROM/XI0/XI2/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM0 XROM/XI0/XI2/NET143 N_WL<4>_XROM/XI0/XI2/MM0_g
+ N_VSS_XROM/XI0/XI2/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM8 N_BL<0>_XROM/XI0/XI1/MM8_d N_WL<3>_XROM/XI0/XI1/MM8_g
+ N_VSS_XROM/XI0/XI1/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM0 XROM/XI0/XI1/NET143 N_WL<2>_XROM/XI0/XI1/MM0_g
+ N_VSS_XROM/XI0/XI1/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM8 N_BL<0>_XROM/XI0/XI0/MM8_d N_WL<1>_XROM/XI0/XI0/MM8_g
+ N_VSS_XROM/XI0/XI0/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM0 XROM/XI0/XI0/NET143 N_WL<0>_XROM/XI0/XI0/MM0_g
+ N_VSS_XROM/XI0/XI0/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM9 XROM/XI1/XI3/NET107 N_WL<15>_XROM/XI1/XI3/MM9_g
+ N_VSS_XROM/XI1/XI3/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM1 N_BL<1>_XROM/XI1/XI3/MM1_d N_WL<14>_XROM/XI1/XI3/MM1_g
+ N_VSS_XROM/XI1/XI3/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM9 XROM/XI1/XI2/NET107 N_WL<13>_XROM/XI1/XI2/MM9_g
+ N_VSS_XROM/XI1/XI2/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM1 N_BL<1>_XROM/XI1/XI2/MM1_d N_WL<12>_XROM/XI1/XI2/MM1_g
+ N_VSS_XROM/XI1/XI2/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM9 XROM/XI1/XI1/NET107 N_WL<11>_XROM/XI1/XI1/MM9_g
+ N_VSS_XROM/XI1/XI1/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM1 N_BL<1>_XROM/XI1/XI1/MM1_d N_WL<10>_XROM/XI1/XI1/MM1_g
+ N_VSS_XROM/XI1/XI1/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM9 XROM/XI1/XI0/NET107 N_WL<9>_XROM/XI1/XI0/MM9_g
+ N_VSS_XROM/XI1/XI0/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM1 N_BL<1>_XROM/XI1/XI0/MM1_d N_WL<8>_XROM/XI1/XI0/MM1_g
+ N_VSS_XROM/XI1/XI0/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM9 XROM/XI0/XI3/NET107 N_WL<7>_XROM/XI0/XI3/MM9_g
+ N_VSS_XROM/XI0/XI3/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM1 N_BL<1>_XROM/XI0/XI3/MM1_d N_WL<6>_XROM/XI0/XI3/MM1_g
+ N_VSS_XROM/XI0/XI3/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM9 XROM/XI0/XI2/NET107 N_WL<5>_XROM/XI0/XI2/MM9_g
+ N_VSS_XROM/XI0/XI2/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM1 N_BL<1>_XROM/XI0/XI2/MM1_d N_WL<4>_XROM/XI0/XI2/MM1_g
+ N_VSS_XROM/XI0/XI2/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM9 XROM/XI0/XI1/NET107 N_WL<3>_XROM/XI0/XI1/MM9_g
+ N_VSS_XROM/XI0/XI1/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM1 N_BL<1>_XROM/XI0/XI1/MM1_d N_WL<2>_XROM/XI0/XI1/MM1_g
+ N_VSS_XROM/XI0/XI1/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM9 XROM/XI0/XI0/NET107 N_WL<1>_XROM/XI0/XI0/MM9_g
+ N_VSS_XROM/XI0/XI0/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM1 N_BL<1>_XROM/XI0/XI0/MM1_d N_WL<0>_XROM/XI0/XI0/MM1_g
+ N_VSS_XROM/XI0/XI0/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM10 N_BL<2>_XROM/XI1/XI3/MM10_d N_WL<15>_XROM/XI1/XI3/MM10_g
+ N_VSS_XROM/XI1/XI3/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM2 XROM/XI1/XI3/NET135 N_WL<14>_XROM/XI1/XI3/MM2_g
+ N_VSS_XROM/XI1/XI3/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM10 N_BL<2>_XROM/XI1/XI2/MM10_d N_WL<13>_XROM/XI1/XI2/MM10_g
+ N_VSS_XROM/XI1/XI2/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM2 XROM/XI1/XI2/NET135 N_WL<12>_XROM/XI1/XI2/MM2_g
+ N_VSS_XROM/XI1/XI2/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM10 N_BL<2>_XROM/XI1/XI1/MM10_d N_WL<11>_XROM/XI1/XI1/MM10_g
+ N_VSS_XROM/XI1/XI1/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM2 XROM/XI1/XI1/NET135 N_WL<10>_XROM/XI1/XI1/MM2_g
+ N_VSS_XROM/XI1/XI1/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM10 N_BL<2>_XROM/XI1/XI0/MM10_d N_WL<9>_XROM/XI1/XI0/MM10_g
+ N_VSS_XROM/XI1/XI0/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM2 XROM/XI1/XI0/NET135 N_WL<8>_XROM/XI1/XI0/MM2_g
+ N_VSS_XROM/XI1/XI0/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM10 N_BL<2>_XROM/XI0/XI3/MM10_d N_WL<7>_XROM/XI0/XI3/MM10_g
+ N_VSS_XROM/XI0/XI3/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM2 XROM/XI0/XI3/NET135 N_WL<6>_XROM/XI0/XI3/MM2_g
+ N_VSS_XROM/XI0/XI3/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM10 N_BL<2>_XROM/XI0/XI2/MM10_d N_WL<5>_XROM/XI0/XI2/MM10_g
+ N_VSS_XROM/XI0/XI2/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM2 XROM/XI0/XI2/NET135 N_WL<4>_XROM/XI0/XI2/MM2_g
+ N_VSS_XROM/XI0/XI2/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM10 N_BL<2>_XROM/XI0/XI1/MM10_d N_WL<3>_XROM/XI0/XI1/MM10_g
+ N_VSS_XROM/XI0/XI1/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM2 XROM/XI0/XI1/NET135 N_WL<2>_XROM/XI0/XI1/MM2_g
+ N_VSS_XROM/XI0/XI1/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM10 N_BL<2>_XROM/XI0/XI0/MM10_d N_WL<1>_XROM/XI0/XI0/MM10_g
+ N_VSS_XROM/XI0/XI0/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM2 XROM/XI0/XI0/NET135 N_WL<0>_XROM/XI0/XI0/MM2_g
+ N_VSS_XROM/XI0/XI0/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM11 XROM/XI1/XI3/NET99 N_WL<15>_XROM/XI1/XI3/MM11_g
+ N_VSS_XROM/XI1/XI3/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM3 N_BL<3>_XROM/XI1/XI3/MM3_d N_WL<14>_XROM/XI1/XI3/MM3_g
+ N_VSS_XROM/XI1/XI3/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM11 XROM/XI1/XI2/NET99 N_WL<13>_XROM/XI1/XI2/MM11_g
+ N_VSS_XROM/XI1/XI2/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM3 N_BL<3>_XROM/XI1/XI2/MM3_d N_WL<12>_XROM/XI1/XI2/MM3_g
+ N_VSS_XROM/XI1/XI2/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM11 XROM/XI1/XI1/NET99 N_WL<11>_XROM/XI1/XI1/MM11_g
+ N_VSS_XROM/XI1/XI1/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM3 N_BL<3>_XROM/XI1/XI1/MM3_d N_WL<10>_XROM/XI1/XI1/MM3_g
+ N_VSS_XROM/XI1/XI1/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM11 XROM/XI1/XI0/NET99 N_WL<9>_XROM/XI1/XI0/MM11_g
+ N_VSS_XROM/XI1/XI0/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM3 N_BL<3>_XROM/XI1/XI0/MM3_d N_WL<8>_XROM/XI1/XI0/MM3_g
+ N_VSS_XROM/XI1/XI0/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM11 XROM/XI0/XI3/NET99 N_WL<7>_XROM/XI0/XI3/MM11_g
+ N_VSS_XROM/XI0/XI3/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM3 N_BL<3>_XROM/XI0/XI3/MM3_d N_WL<6>_XROM/XI0/XI3/MM3_g
+ N_VSS_XROM/XI0/XI3/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM11 XROM/XI0/XI2/NET99 N_WL<5>_XROM/XI0/XI2/MM11_g
+ N_VSS_XROM/XI0/XI2/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM3 N_BL<3>_XROM/XI0/XI2/MM3_d N_WL<4>_XROM/XI0/XI2/MM3_g
+ N_VSS_XROM/XI0/XI2/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM11 XROM/XI0/XI1/NET99 N_WL<3>_XROM/XI0/XI1/MM11_g
+ N_VSS_XROM/XI0/XI1/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM3 N_BL<3>_XROM/XI0/XI1/MM3_d N_WL<2>_XROM/XI0/XI1/MM3_g
+ N_VSS_XROM/XI0/XI1/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM11 XROM/XI0/XI0/NET99 N_WL<1>_XROM/XI0/XI0/MM11_g
+ N_VSS_XROM/XI0/XI0/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM3 N_BL<3>_XROM/XI0/XI0/MM3_d N_WL<0>_XROM/XI0/XI0/MM3_g
+ N_VSS_XROM/XI0/XI0/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM12 N_BL<4>_XROM/XI1/XI3/MM12_d N_WL<15>_XROM/XI1/XI3/MM12_g
+ N_VSS_XROM/XI1/XI3/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM4 XROM/XI1/XI3/NET127 N_WL<14>_XROM/XI1/XI3/MM4_g
+ N_VSS_XROM/XI1/XI3/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM12 N_BL<4>_XROM/XI1/XI2/MM12_d N_WL<13>_XROM/XI1/XI2/MM12_g
+ N_VSS_XROM/XI1/XI2/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM4 XROM/XI1/XI2/NET127 N_WL<12>_XROM/XI1/XI2/MM4_g
+ N_VSS_XROM/XI1/XI2/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM12 N_BL<4>_XROM/XI1/XI1/MM12_d N_WL<11>_XROM/XI1/XI1/MM12_g
+ N_VSS_XROM/XI1/XI1/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM4 XROM/XI1/XI1/NET127 N_WL<10>_XROM/XI1/XI1/MM4_g
+ N_VSS_XROM/XI1/XI1/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM12 N_BL<4>_XROM/XI1/XI0/MM12_d N_WL<9>_XROM/XI1/XI0/MM12_g
+ N_VSS_XROM/XI1/XI0/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM4 XROM/XI1/XI0/NET127 N_WL<8>_XROM/XI1/XI0/MM4_g
+ N_VSS_XROM/XI1/XI0/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM12 N_BL<4>_XROM/XI0/XI3/MM12_d N_WL<7>_XROM/XI0/XI3/MM12_g
+ N_VSS_XROM/XI0/XI3/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM4 XROM/XI0/XI3/NET127 N_WL<6>_XROM/XI0/XI3/MM4_g
+ N_VSS_XROM/XI0/XI3/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM12 N_BL<4>_XROM/XI0/XI2/MM12_d N_WL<5>_XROM/XI0/XI2/MM12_g
+ N_VSS_XROM/XI0/XI2/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM4 XROM/XI0/XI2/NET127 N_WL<4>_XROM/XI0/XI2/MM4_g
+ N_VSS_XROM/XI0/XI2/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM12 N_BL<4>_XROM/XI0/XI1/MM12_d N_WL<3>_XROM/XI0/XI1/MM12_g
+ N_VSS_XROM/XI0/XI1/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM4 XROM/XI0/XI1/NET127 N_WL<2>_XROM/XI0/XI1/MM4_g
+ N_VSS_XROM/XI0/XI1/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM12 N_BL<4>_XROM/XI0/XI0/MM12_d N_WL<1>_XROM/XI0/XI0/MM12_g
+ N_VSS_XROM/XI0/XI0/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM4 XROM/XI0/XI0/NET127 N_WL<0>_XROM/XI0/XI0/MM4_g
+ N_VSS_XROM/XI0/XI0/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM13 XROM/XI1/XI3/NET91 N_WL<15>_XROM/XI1/XI3/MM13_g
+ N_VSS_XROM/XI1/XI3/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM5 N_BL<5>_XROM/XI1/XI3/MM5_d N_WL<14>_XROM/XI1/XI3/MM5_g
+ N_VSS_XROM/XI1/XI3/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM13 XROM/XI1/XI2/NET91 N_WL<13>_XROM/XI1/XI2/MM13_g
+ N_VSS_XROM/XI1/XI2/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM5 N_BL<5>_XROM/XI1/XI2/MM5_d N_WL<12>_XROM/XI1/XI2/MM5_g
+ N_VSS_XROM/XI1/XI2/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM13 XROM/XI1/XI1/NET91 N_WL<11>_XROM/XI1/XI1/MM13_g
+ N_VSS_XROM/XI1/XI1/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM5 N_BL<5>_XROM/XI1/XI1/MM5_d N_WL<10>_XROM/XI1/XI1/MM5_g
+ N_VSS_XROM/XI1/XI1/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM13 XROM/XI1/XI0/NET91 N_WL<9>_XROM/XI1/XI0/MM13_g
+ N_VSS_XROM/XI1/XI0/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM5 N_BL<5>_XROM/XI1/XI0/MM5_d N_WL<8>_XROM/XI1/XI0/MM5_g
+ N_VSS_XROM/XI1/XI0/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM13 XROM/XI0/XI3/NET91 N_WL<7>_XROM/XI0/XI3/MM13_g
+ N_VSS_XROM/XI0/XI3/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM5 N_BL<5>_XROM/XI0/XI3/MM5_d N_WL<6>_XROM/XI0/XI3/MM5_g
+ N_VSS_XROM/XI0/XI3/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM13 XROM/XI0/XI2/NET91 N_WL<5>_XROM/XI0/XI2/MM13_g
+ N_VSS_XROM/XI0/XI2/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM5 N_BL<5>_XROM/XI0/XI2/MM5_d N_WL<4>_XROM/XI0/XI2/MM5_g
+ N_VSS_XROM/XI0/XI2/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM13 XROM/XI0/XI1/NET91 N_WL<3>_XROM/XI0/XI1/MM13_g
+ N_VSS_XROM/XI0/XI1/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM5 N_BL<5>_XROM/XI0/XI1/MM5_d N_WL<2>_XROM/XI0/XI1/MM5_g
+ N_VSS_XROM/XI0/XI1/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM13 XROM/XI0/XI0/NET91 N_WL<1>_XROM/XI0/XI0/MM13_g
+ N_VSS_XROM/XI0/XI0/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM5 N_BL<5>_XROM/XI0/XI0/MM5_d N_WL<0>_XROM/XI0/XI0/MM5_g
+ N_VSS_XROM/XI0/XI0/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM14 N_BL<6>_XROM/XI1/XI3/MM14_d N_WL<15>_XROM/XI1/XI3/MM14_g
+ N_VSS_XROM/XI1/XI3/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM6 XROM/XI1/XI3/NET119 N_WL<14>_XROM/XI1/XI3/MM6_g
+ N_VSS_XROM/XI1/XI3/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM14 N_BL<6>_XROM/XI1/XI2/MM14_d N_WL<13>_XROM/XI1/XI2/MM14_g
+ N_VSS_XROM/XI1/XI2/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM6 XROM/XI1/XI2/NET119 N_WL<12>_XROM/XI1/XI2/MM6_g
+ N_VSS_XROM/XI1/XI2/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM14 N_BL<6>_XROM/XI1/XI1/MM14_d N_WL<11>_XROM/XI1/XI1/MM14_g
+ N_VSS_XROM/XI1/XI1/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM6 XROM/XI1/XI1/NET119 N_WL<10>_XROM/XI1/XI1/MM6_g
+ N_VSS_XROM/XI1/XI1/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM14 N_BL<6>_XROM/XI1/XI0/MM14_d N_WL<9>_XROM/XI1/XI0/MM14_g
+ N_VSS_XROM/XI1/XI0/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM6 XROM/XI1/XI0/NET119 N_WL<8>_XROM/XI1/XI0/MM6_g
+ N_VSS_XROM/XI1/XI0/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM14 N_BL<6>_XROM/XI0/XI3/MM14_d N_WL<7>_XROM/XI0/XI3/MM14_g
+ N_VSS_XROM/XI0/XI3/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM6 XROM/XI0/XI3/NET119 N_WL<6>_XROM/XI0/XI3/MM6_g
+ N_VSS_XROM/XI0/XI3/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM14 N_BL<6>_XROM/XI0/XI2/MM14_d N_WL<5>_XROM/XI0/XI2/MM14_g
+ N_VSS_XROM/XI0/XI2/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM6 XROM/XI0/XI2/NET119 N_WL<4>_XROM/XI0/XI2/MM6_g
+ N_VSS_XROM/XI0/XI2/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM14 N_BL<6>_XROM/XI0/XI1/MM14_d N_WL<3>_XROM/XI0/XI1/MM14_g
+ N_VSS_XROM/XI0/XI1/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM6 XROM/XI0/XI1/NET119 N_WL<2>_XROM/XI0/XI1/MM6_g
+ N_VSS_XROM/XI0/XI1/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM14 N_BL<6>_XROM/XI0/XI0/MM14_d N_WL<1>_XROM/XI0/XI0/MM14_g
+ N_VSS_XROM/XI0/XI0/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM6 XROM/XI0/XI0/NET119 N_WL<0>_XROM/XI0/XI0/MM6_g
+ N_VSS_XROM/XI0/XI0/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM15 XROM/XI1/XI3/NET83 N_WL<15>_XROM/XI1/XI3/MM15_g
+ N_VSS_XROM/XI1/XI3/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI3/MM7 N_BL<7>_XROM/XI1/XI3/MM7_d N_WL<14>_XROM/XI1/XI3/MM7_g
+ N_VSS_XROM/XI1/XI3/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM15 XROM/XI1/XI2/NET83 N_WL<13>_XROM/XI1/XI2/MM15_g
+ N_VSS_XROM/XI1/XI2/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI2/MM7 N_BL<7>_XROM/XI1/XI2/MM7_d N_WL<12>_XROM/XI1/XI2/MM7_g
+ N_VSS_XROM/XI1/XI2/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM15 XROM/XI1/XI1/NET83 N_WL<11>_XROM/XI1/XI1/MM15_g
+ N_VSS_XROM/XI1/XI1/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI1/MM7 N_BL<7>_XROM/XI1/XI1/MM7_d N_WL<10>_XROM/XI1/XI1/MM7_g
+ N_VSS_XROM/XI1/XI1/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM15 XROM/XI1/XI0/NET83 N_WL<9>_XROM/XI1/XI0/MM15_g
+ N_VSS_XROM/XI1/XI0/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI0/MM7 N_BL<7>_XROM/XI1/XI0/MM7_d N_WL<8>_XROM/XI1/XI0/MM7_g
+ N_VSS_XROM/XI1/XI0/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM15 XROM/XI0/XI3/NET83 N_WL<7>_XROM/XI0/XI3/MM15_g
+ N_VSS_XROM/XI0/XI3/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI3/MM7 N_BL<7>_XROM/XI0/XI3/MM7_d N_WL<6>_XROM/XI0/XI3/MM7_g
+ N_VSS_XROM/XI0/XI3/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM15 XROM/XI0/XI2/NET83 N_WL<5>_XROM/XI0/XI2/MM15_g
+ N_VSS_XROM/XI0/XI2/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI2/MM7 N_BL<7>_XROM/XI0/XI2/MM7_d N_WL<4>_XROM/XI0/XI2/MM7_g
+ N_VSS_XROM/XI0/XI2/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM15 XROM/XI0/XI1/NET83 N_WL<3>_XROM/XI0/XI1/MM15_g
+ N_VSS_XROM/XI0/XI1/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI1/MM7 N_BL<7>_XROM/XI0/XI1/MM7_d N_WL<2>_XROM/XI0/XI1/MM7_g
+ N_VSS_XROM/XI0/XI1/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM15 XROM/XI0/XI0/NET83 N_WL<1>_XROM/XI0/XI0/MM15_g
+ N_VSS_XROM/XI0/XI0/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI0/MM7 N_BL<7>_XROM/XI0/XI0/MM7_d N_WL<0>_XROM/XI0/XI0/MM7_g
+ N_VSS_XROM/XI0/XI0/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM8 N_BL<8>_XROM/XI1/XI7/MM8_d N_WL<15>_XROM/XI1/XI7/MM8_g
+ N_VSS_XROM/XI1/XI7/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM0 XROM/XI1/XI7/NET143 N_WL<14>_XROM/XI1/XI7/MM0_g
+ N_VSS_XROM/XI1/XI7/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM8 N_BL<8>_XROM/XI1/XI6/MM8_d N_WL<13>_XROM/XI1/XI6/MM8_g
+ N_VSS_XROM/XI1/XI6/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM0 XROM/XI1/XI6/NET143 N_WL<12>_XROM/XI1/XI6/MM0_g
+ N_VSS_XROM/XI1/XI6/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM8 N_BL<8>_XROM/XI1/XI5/MM8_d N_WL<11>_XROM/XI1/XI5/MM8_g
+ N_VSS_XROM/XI1/XI5/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM0 XROM/XI1/XI5/NET143 N_WL<10>_XROM/XI1/XI5/MM0_g
+ N_VSS_XROM/XI1/XI5/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM8 N_BL<8>_XROM/XI1/XI4/MM8_d N_WL<9>_XROM/XI1/XI4/MM8_g
+ N_VSS_XROM/XI1/XI4/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM0 XROM/XI1/XI4/NET143 N_WL<8>_XROM/XI1/XI4/MM0_g
+ N_VSS_XROM/XI1/XI4/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM8 N_BL<8>_XROM/XI0/XI7/MM8_d N_WL<7>_XROM/XI0/XI7/MM8_g
+ N_VSS_XROM/XI0/XI7/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM0 XROM/XI0/XI7/NET143 N_WL<6>_XROM/XI0/XI7/MM0_g
+ N_VSS_XROM/XI0/XI7/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM8 N_BL<8>_XROM/XI0/XI6/MM8_d N_WL<5>_XROM/XI0/XI6/MM8_g
+ N_VSS_XROM/XI0/XI6/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM0 XROM/XI0/XI6/NET143 N_WL<4>_XROM/XI0/XI6/MM0_g
+ N_VSS_XROM/XI0/XI6/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM8 N_BL<8>_XROM/XI0/XI5/MM8_d N_WL<3>_XROM/XI0/XI5/MM8_g
+ N_VSS_XROM/XI0/XI5/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM0 XROM/XI0/XI5/NET143 N_WL<2>_XROM/XI0/XI5/MM0_g
+ N_VSS_XROM/XI0/XI5/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM8 N_BL<8>_XROM/XI0/XI4/MM8_d N_WL<1>_XROM/XI0/XI4/MM8_g
+ N_VSS_XROM/XI0/XI4/MM8_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM0 XROM/XI0/XI4/NET143 N_WL<0>_XROM/XI0/XI4/MM0_g
+ N_VSS_XROM/XI0/XI4/MM0_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM9 XROM/XI1/XI7/NET107 N_WL<15>_XROM/XI1/XI7/MM9_g
+ N_VSS_XROM/XI1/XI7/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM1 N_BL<9>_XROM/XI1/XI7/MM1_d N_WL<14>_XROM/XI1/XI7/MM1_g
+ N_VSS_XROM/XI1/XI7/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM9 XROM/XI1/XI6/NET107 N_WL<13>_XROM/XI1/XI6/MM9_g
+ N_VSS_XROM/XI1/XI6/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM1 N_BL<9>_XROM/XI1/XI6/MM1_d N_WL<12>_XROM/XI1/XI6/MM1_g
+ N_VSS_XROM/XI1/XI6/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM9 XROM/XI1/XI5/NET107 N_WL<11>_XROM/XI1/XI5/MM9_g
+ N_VSS_XROM/XI1/XI5/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM1 N_BL<9>_XROM/XI1/XI5/MM1_d N_WL<10>_XROM/XI1/XI5/MM1_g
+ N_VSS_XROM/XI1/XI5/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM9 XROM/XI1/XI4/NET107 N_WL<9>_XROM/XI1/XI4/MM9_g
+ N_VSS_XROM/XI1/XI4/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM1 N_BL<9>_XROM/XI1/XI4/MM1_d N_WL<8>_XROM/XI1/XI4/MM1_g
+ N_VSS_XROM/XI1/XI4/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM9 XROM/XI0/XI7/NET107 N_WL<7>_XROM/XI0/XI7/MM9_g
+ N_VSS_XROM/XI0/XI7/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM1 N_BL<9>_XROM/XI0/XI7/MM1_d N_WL<6>_XROM/XI0/XI7/MM1_g
+ N_VSS_XROM/XI0/XI7/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM9 XROM/XI0/XI6/NET107 N_WL<5>_XROM/XI0/XI6/MM9_g
+ N_VSS_XROM/XI0/XI6/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM1 N_BL<9>_XROM/XI0/XI6/MM1_d N_WL<4>_XROM/XI0/XI6/MM1_g
+ N_VSS_XROM/XI0/XI6/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM9 XROM/XI0/XI5/NET107 N_WL<3>_XROM/XI0/XI5/MM9_g
+ N_VSS_XROM/XI0/XI5/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM1 N_BL<9>_XROM/XI0/XI5/MM1_d N_WL<2>_XROM/XI0/XI5/MM1_g
+ N_VSS_XROM/XI0/XI5/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM9 XROM/XI0/XI4/NET107 N_WL<1>_XROM/XI0/XI4/MM9_g
+ N_VSS_XROM/XI0/XI4/MM9_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM1 N_BL<9>_XROM/XI0/XI4/MM1_d N_WL<0>_XROM/XI0/XI4/MM1_g
+ N_VSS_XROM/XI0/XI4/MM1_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM10 N_BL<10>_XROM/XI1/XI7/MM10_d N_WL<15>_XROM/XI1/XI7/MM10_g
+ N_VSS_XROM/XI1/XI7/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM2 XROM/XI1/XI7/NET135 N_WL<14>_XROM/XI1/XI7/MM2_g
+ N_VSS_XROM/XI1/XI7/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM10 N_BL<10>_XROM/XI1/XI6/MM10_d N_WL<13>_XROM/XI1/XI6/MM10_g
+ N_VSS_XROM/XI1/XI6/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM2 XROM/XI1/XI6/NET135 N_WL<12>_XROM/XI1/XI6/MM2_g
+ N_VSS_XROM/XI1/XI6/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM10 N_BL<10>_XROM/XI1/XI5/MM10_d N_WL<11>_XROM/XI1/XI5/MM10_g
+ N_VSS_XROM/XI1/XI5/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM2 XROM/XI1/XI5/NET135 N_WL<10>_XROM/XI1/XI5/MM2_g
+ N_VSS_XROM/XI1/XI5/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM10 N_BL<10>_XROM/XI1/XI4/MM10_d N_WL<9>_XROM/XI1/XI4/MM10_g
+ N_VSS_XROM/XI1/XI4/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM2 XROM/XI1/XI4/NET135 N_WL<8>_XROM/XI1/XI4/MM2_g
+ N_VSS_XROM/XI1/XI4/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM10 N_BL<10>_XROM/XI0/XI7/MM10_d N_WL<7>_XROM/XI0/XI7/MM10_g
+ N_VSS_XROM/XI0/XI7/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM2 XROM/XI0/XI7/NET135 N_WL<6>_XROM/XI0/XI7/MM2_g
+ N_VSS_XROM/XI0/XI7/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM10 N_BL<10>_XROM/XI0/XI6/MM10_d N_WL<5>_XROM/XI0/XI6/MM10_g
+ N_VSS_XROM/XI0/XI6/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM2 XROM/XI0/XI6/NET135 N_WL<4>_XROM/XI0/XI6/MM2_g
+ N_VSS_XROM/XI0/XI6/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM10 N_BL<10>_XROM/XI0/XI5/MM10_d N_WL<3>_XROM/XI0/XI5/MM10_g
+ N_VSS_XROM/XI0/XI5/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM2 XROM/XI0/XI5/NET135 N_WL<2>_XROM/XI0/XI5/MM2_g
+ N_VSS_XROM/XI0/XI5/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM10 N_BL<10>_XROM/XI0/XI4/MM10_d N_WL<1>_XROM/XI0/XI4/MM10_g
+ N_VSS_XROM/XI0/XI4/MM10_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM2 XROM/XI0/XI4/NET135 N_WL<0>_XROM/XI0/XI4/MM2_g
+ N_VSS_XROM/XI0/XI4/MM2_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM11 XROM/XI1/XI7/NET99 N_WL<15>_XROM/XI1/XI7/MM11_g
+ N_VSS_XROM/XI1/XI7/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM3 N_BL<11>_XROM/XI1/XI7/MM3_d N_WL<14>_XROM/XI1/XI7/MM3_g
+ N_VSS_XROM/XI1/XI7/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM11 XROM/XI1/XI6/NET99 N_WL<13>_XROM/XI1/XI6/MM11_g
+ N_VSS_XROM/XI1/XI6/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM3 N_BL<11>_XROM/XI1/XI6/MM3_d N_WL<12>_XROM/XI1/XI6/MM3_g
+ N_VSS_XROM/XI1/XI6/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM11 XROM/XI1/XI5/NET99 N_WL<11>_XROM/XI1/XI5/MM11_g
+ N_VSS_XROM/XI1/XI5/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM3 N_BL<11>_XROM/XI1/XI5/MM3_d N_WL<10>_XROM/XI1/XI5/MM3_g
+ N_VSS_XROM/XI1/XI5/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM11 XROM/XI1/XI4/NET99 N_WL<9>_XROM/XI1/XI4/MM11_g
+ N_VSS_XROM/XI1/XI4/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM3 N_BL<11>_XROM/XI1/XI4/MM3_d N_WL<8>_XROM/XI1/XI4/MM3_g
+ N_VSS_XROM/XI1/XI4/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM11 XROM/XI0/XI7/NET99 N_WL<7>_XROM/XI0/XI7/MM11_g
+ N_VSS_XROM/XI0/XI7/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM3 N_BL<11>_XROM/XI0/XI7/MM3_d N_WL<6>_XROM/XI0/XI7/MM3_g
+ N_VSS_XROM/XI0/XI7/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM13 XROM/XI0/XI6/NET91 N_WL<5>_XROM/XI0/XI6/MM13_g
+ N_VSS_XROM/XI0/XI6/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM3 N_BL<11>_XROM/XI0/XI6/MM3_d N_WL<4>_XROM/XI0/XI6/MM3_g
+ N_VSS_XROM/XI0/XI6/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM13 XROM/XI0/XI5/NET91 N_WL<3>_XROM/XI0/XI5/MM13_g
+ N_VSS_XROM/XI0/XI5/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM3 N_BL<11>_XROM/XI0/XI5/MM3_d N_WL<2>_XROM/XI0/XI5/MM3_g
+ N_VSS_XROM/XI0/XI5/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM13 XROM/XI0/XI4/NET91 N_WL<1>_XROM/XI0/XI4/MM13_g
+ N_VSS_XROM/XI0/XI4/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM3 N_BL<11>_XROM/XI0/XI4/MM3_d N_WL<0>_XROM/XI0/XI4/MM3_g
+ N_VSS_XROM/XI0/XI4/MM3_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM12 N_BL<12>_XROM/XI1/XI7/MM12_d N_WL<15>_XROM/XI1/XI7/MM12_g
+ N_VSS_XROM/XI1/XI7/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM4 XROM/XI1/XI7/NET127 N_WL<14>_XROM/XI1/XI7/MM4_g
+ N_VSS_XROM/XI1/XI7/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM12 N_BL<12>_XROM/XI1/XI6/MM12_d N_WL<13>_XROM/XI1/XI6/MM12_g
+ N_VSS_XROM/XI1/XI6/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM4 XROM/XI1/XI6/NET127 N_WL<12>_XROM/XI1/XI6/MM4_g
+ N_VSS_XROM/XI1/XI6/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM12 N_BL<12>_XROM/XI1/XI5/MM12_d N_WL<11>_XROM/XI1/XI5/MM12_g
+ N_VSS_XROM/XI1/XI5/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM4 XROM/XI1/XI5/NET127 N_WL<10>_XROM/XI1/XI5/MM4_g
+ N_VSS_XROM/XI1/XI5/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM12 N_BL<12>_XROM/XI1/XI4/MM12_d N_WL<9>_XROM/XI1/XI4/MM12_g
+ N_VSS_XROM/XI1/XI4/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM4 XROM/XI1/XI4/NET127 N_WL<8>_XROM/XI1/XI4/MM4_g
+ N_VSS_XROM/XI1/XI4/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM12 N_BL<12>_XROM/XI0/XI7/MM12_d N_WL<7>_XROM/XI0/XI7/MM12_g
+ N_VSS_XROM/XI0/XI7/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM4 XROM/XI0/XI7/NET127 N_WL<6>_XROM/XI0/XI7/MM4_g
+ N_VSS_XROM/XI0/XI7/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM12 N_BL<12>_XROM/XI0/XI6/MM12_d N_WL<5>_XROM/XI0/XI6/MM12_g
+ N_VSS_XROM/XI0/XI6/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM6 XROM/XI0/XI6/NET119 N_WL<4>_XROM/XI0/XI6/MM6_g
+ N_VSS_XROM/XI0/XI6/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM12 N_BL<12>_XROM/XI0/XI5/MM12_d N_WL<3>_XROM/XI0/XI5/MM12_g
+ N_VSS_XROM/XI0/XI5/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM6 XROM/XI0/XI5/NET119 N_WL<2>_XROM/XI0/XI5/MM6_g
+ N_VSS_XROM/XI0/XI5/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM12 N_BL<12>_XROM/XI0/XI4/MM12_d N_WL<1>_XROM/XI0/XI4/MM12_g
+ N_VSS_XROM/XI0/XI4/MM12_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM6 XROM/XI0/XI4/NET119 N_WL<0>_XROM/XI0/XI4/MM6_g
+ N_VSS_XROM/XI0/XI4/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM15 XROM/XI1/XI7/NET83 N_WL<15>_XROM/XI1/XI7/MM15_g
+ N_VSS_XROM/XI1/XI7/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM5 N_BL<13>_XROM/XI1/XI7/MM5_d N_WL<14>_XROM/XI1/XI7/MM5_g
+ N_VSS_XROM/XI1/XI7/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM15 XROM/XI1/XI6/NET83 N_WL<13>_XROM/XI1/XI6/MM15_g
+ N_VSS_XROM/XI1/XI6/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM5 N_BL<13>_XROM/XI1/XI6/MM5_d N_WL<12>_XROM/XI1/XI6/MM5_g
+ N_VSS_XROM/XI1/XI6/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM15 XROM/XI1/XI5/NET83 N_WL<11>_XROM/XI1/XI5/MM15_g
+ N_VSS_XROM/XI1/XI5/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM5 N_BL<13>_XROM/XI1/XI5/MM5_d N_WL<10>_XROM/XI1/XI5/MM5_g
+ N_VSS_XROM/XI1/XI5/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM15 XROM/XI1/XI4/NET83 N_WL<9>_XROM/XI1/XI4/MM15_g
+ N_VSS_XROM/XI1/XI4/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM5 N_BL<13>_XROM/XI1/XI4/MM5_d N_WL<8>_XROM/XI1/XI4/MM5_g
+ N_VSS_XROM/XI1/XI4/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM15 XROM/XI0/XI7/NET83 N_WL<7>_XROM/XI0/XI7/MM15_g
+ N_VSS_XROM/XI0/XI7/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM5 N_BL<13>_XROM/XI0/XI7/MM5_d N_WL<6>_XROM/XI0/XI7/MM5_g
+ N_VSS_XROM/XI0/XI7/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM15 XROM/XI0/XI6/NET83 N_WL<5>_XROM/XI0/XI6/MM15_g
+ N_VSS_XROM/XI0/XI6/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM5 N_BL<13>_XROM/XI0/XI6/MM5_d N_WL<4>_XROM/XI0/XI6/MM5_g
+ N_VSS_XROM/XI0/XI6/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM15 XROM/XI0/XI5/NET83 N_WL<3>_XROM/XI0/XI5/MM15_g
+ N_VSS_XROM/XI0/XI5/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM5 N_BL<13>_XROM/XI0/XI5/MM5_d N_WL<2>_XROM/XI0/XI5/MM5_g
+ N_VSS_XROM/XI0/XI5/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM15 XROM/XI0/XI4/NET83 N_WL<1>_XROM/XI0/XI4/MM15_g
+ N_VSS_XROM/XI0/XI4/MM15_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM5 N_BL<13>_XROM/XI0/XI4/MM5_d N_WL<0>_XROM/XI0/XI4/MM5_g
+ N_VSS_XROM/XI0/XI4/MM5_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM14 N_BL<14>_XROM/XI1/XI7/MM14_d N_WL<15>_XROM/XI1/XI7/MM14_g
+ N_VSS_XROM/XI1/XI7/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM6 XROM/XI1/XI7/NET119 N_WL<14>_XROM/XI1/XI7/MM6_g
+ N_VSS_XROM/XI1/XI7/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM14 N_BL<14>_XROM/XI1/XI6/MM14_d N_WL<13>_XROM/XI1/XI6/MM14_g
+ N_VSS_XROM/XI1/XI6/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM6 XROM/XI1/XI6/NET119 N_WL<12>_XROM/XI1/XI6/MM6_g
+ N_VSS_XROM/XI1/XI6/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM14 N_BL<14>_XROM/XI1/XI5/MM14_d N_WL<11>_XROM/XI1/XI5/MM14_g
+ N_VSS_XROM/XI1/XI5/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM6 XROM/XI1/XI5/NET119 N_WL<10>_XROM/XI1/XI5/MM6_g
+ N_VSS_XROM/XI1/XI5/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM14 N_BL<14>_XROM/XI1/XI4/MM14_d N_WL<9>_XROM/XI1/XI4/MM14_g
+ N_VSS_XROM/XI1/XI4/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM6 XROM/XI1/XI4/NET119 N_WL<8>_XROM/XI1/XI4/MM6_g
+ N_VSS_XROM/XI1/XI4/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM14 N_BL<14>_XROM/XI0/XI7/MM14_d N_WL<7>_XROM/XI0/XI7/MM14_g
+ N_VSS_XROM/XI0/XI7/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM6 XROM/XI0/XI7/NET119 N_WL<6>_XROM/XI0/XI7/MM6_g
+ N_VSS_XROM/XI0/XI7/MM6_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM14 N_BL<14>_XROM/XI0/XI6/MM14_d N_WL<5>_XROM/XI0/XI6/MM14_g
+ N_VSS_XROM/XI0/XI6/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM4 XROM/XI0/XI6/NET127 N_WL<4>_XROM/XI0/XI6/MM4_g
+ N_VSS_XROM/XI0/XI6/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM14 N_BL<14>_XROM/XI0/XI5/MM14_d N_WL<3>_XROM/XI0/XI5/MM14_g
+ N_VSS_XROM/XI0/XI5/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM4 XROM/XI0/XI5/NET127 N_WL<2>_XROM/XI0/XI5/MM4_g
+ N_VSS_XROM/XI0/XI5/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM14 N_BL<14>_XROM/XI0/XI4/MM14_d N_WL<1>_XROM/XI0/XI4/MM14_g
+ N_VSS_XROM/XI0/XI4/MM14_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM4 XROM/XI0/XI4/NET127 N_WL<0>_XROM/XI0/XI4/MM4_g
+ N_VSS_XROM/XI0/XI4/MM4_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM13 XROM/XI1/XI7/NET91 N_WL<15>_XROM/XI1/XI7/MM13_g
+ N_VSS_XROM/XI1/XI7/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI7/MM7 N_BL<15>_XROM/XI1/XI7/MM7_d N_WL<14>_XROM/XI1/XI7/MM7_g
+ N_VSS_XROM/XI1/XI7/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM13 XROM/XI1/XI6/NET91 N_WL<13>_XROM/XI1/XI6/MM13_g
+ N_VSS_XROM/XI1/XI6/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI6/MM7 N_BL<15>_XROM/XI1/XI6/MM7_d N_WL<12>_XROM/XI1/XI6/MM7_g
+ N_VSS_XROM/XI1/XI6/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM13 XROM/XI1/XI5/NET91 N_WL<11>_XROM/XI1/XI5/MM13_g
+ N_VSS_XROM/XI1/XI5/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI5/MM7 N_BL<15>_XROM/XI1/XI5/MM7_d N_WL<10>_XROM/XI1/XI5/MM7_g
+ N_VSS_XROM/XI1/XI5/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM13 XROM/XI1/XI4/NET91 N_WL<9>_XROM/XI1/XI4/MM13_g
+ N_VSS_XROM/XI1/XI4/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI1/XI4/MM7 N_BL<15>_XROM/XI1/XI4/MM7_d N_WL<8>_XROM/XI1/XI4/MM7_g
+ N_VSS_XROM/XI1/XI4/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM13 XROM/XI0/XI7/NET91 N_WL<7>_XROM/XI0/XI7/MM13_g
+ N_VSS_XROM/XI0/XI7/MM13_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI7/MM7 N_BL<15>_XROM/XI0/XI7/MM7_d N_WL<6>_XROM/XI0/XI7/MM7_g
+ N_VSS_XROM/XI0/XI7/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM11 XROM/XI0/XI6/NET99 N_WL<5>_XROM/XI0/XI6/MM11_g
+ N_VSS_XROM/XI0/XI6/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI6/MM7 N_BL<15>_XROM/XI0/XI6/MM7_d N_WL<4>_XROM/XI0/XI6/MM7_g
+ N_VSS_XROM/XI0/XI6/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM11 XROM/XI0/XI5/NET99 N_WL<3>_XROM/XI0/XI5/MM11_g
+ N_VSS_XROM/XI0/XI5/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI5/MM7 N_BL<15>_XROM/XI0/XI5/MM7_d N_WL<2>_XROM/XI0/XI5/MM7_g
+ N_VSS_XROM/XI0/XI5/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM11 XROM/XI0/XI4/NET99 N_WL<1>_XROM/XI0/XI4/MM11_g
+ N_VSS_XROM/XI0/XI4/MM11_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXROM/XI0/XI4/MM7 N_BL<15>_XROM/XI0/XI4/MM7_d N_WL<0>_XROM/XI0/XI4/MM7_g
+ N_VSS_XROM/XI0/XI4/MM7_s N_VSS_XDFF_Timing_control/XI3/MM0_b N_18 L=1.8e-07
+ W=4.7e-07 AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
c_1 XROM/XI7/XI3/NET119 0 0.14368f
c_2 XROM/XI7/XI3/NET107 0 0.180473f
c_3 XROM/XI7/XI7/NET135 0 0.176433f
c_4 XROM/XI7/XI3/NET99 0 0.180473f
c_5 XROM/XI7/XI3/NET135 0 0.176433f
c_6 XROM/XI7/XI3/NET91 0 0.180473f
c_7 XROM/XI7/XI7/NET119 0 0.176433f
c_8 XROM/XI7/XI3/NET83 0 0.180502f
c_9 XROM/XI7/XI3/NET127 0 0.176433f
c_10 XROM/XI7/XI7/NET107 0 0.180475f
c_11 XROM/XI7/XI7/NET127 0 0.176433f
c_12 XROM/XI7/XI7/NET99 0 0.180473f
c_13 XROM/XI7/XI7/NET143 0 0.176433f
c_14 XROM/XI7/XI7/NET91 0 0.180473f
c_15 XROM/XI7/XI3/NET143 0 0.176433f
c_16 XROM/XI7/XI7/NET83 0 0.137954f
c_17 XROM/XI7/XI2/NET143 0 0.138821f
c_18 XROM/XI7/XI2/NET107 0 0.176433f
c_19 XROM/XI7/XI2/NET135 0 0.176433f
c_20 XROM/XI7/XI2/NET99 0 0.176433f
c_21 XROM/XI7/XI2/NET127 0 0.176433f
c_22 XROM/XI7/XI2/NET91 0 0.176433f
c_23 XROM/XI7/XI2/NET119 0 0.176433f
c_24 XROM/XI7/XI2/NET83 0 0.176433f
c_25 XROM/XI7/XI6/NET143 0 0.176433f
c_26 XROM/XI7/XI6/NET107 0 0.176433f
c_27 XROM/XI7/XI6/NET135 0 0.176433f
c_28 XROM/XI7/XI6/NET99 0 0.176433f
c_29 XROM/XI7/XI6/NET127 0 0.176433f
c_30 XROM/XI7/XI6/NET91 0 0.176433f
c_31 XROM/XI7/XI6/NET119 0 0.176433f
c_32 XROM/XI7/XI6/NET83 0 0.136314f
c_33 XROM/XI7/XI1/NET143 0 0.142339f
c_34 XROM/XI7/XI1/NET107 0 0.176433f
c_35 XROM/XI7/XI1/NET135 0 0.176433f
c_36 XROM/XI7/XI1/NET99 0 0.176433f
c_37 XROM/XI7/XI1/NET127 0 0.176433f
c_38 XROM/XI7/XI1/NET91 0 0.176433f
c_39 XROM/XI7/XI1/NET119 0 0.176433f
c_40 XROM/XI7/XI1/NET83 0 0.176433f
c_41 XROM/XI7/XI5/NET143 0 0.176433f
c_42 XROM/XI7/XI5/NET107 0 0.176433f
c_43 XROM/XI7/XI5/NET135 0 0.176433f
c_44 XROM/XI7/XI5/NET99 0 0.176433f
c_45 XROM/XI7/XI5/NET127 0 0.176433f
c_46 XROM/XI7/XI5/NET91 0 0.176433f
c_47 XROM/XI7/XI5/NET119 0 0.176433f
c_48 XROM/XI7/XI5/NET83 0 0.136314f
c_49 XROM/XI7/XI0/NET143 0 0.14368f
c_50 XROM/XI7/XI0/NET107 0 0.176433f
c_51 XROM/XI7/XI0/NET135 0 0.176433f
c_52 XROM/XI7/XI0/NET99 0 0.176433f
c_53 XROM/XI7/XI0/NET127 0 0.176433f
c_54 XROM/XI7/XI0/NET91 0 0.176433f
c_55 XROM/XI7/XI0/NET119 0 0.176433f
c_56 XROM/XI7/XI0/NET83 0 0.176433f
c_57 XROM/XI7/XI4/NET143 0 0.176433f
c_58 XROM/XI7/XI4/NET107 0 0.176433f
c_59 XROM/XI7/XI4/NET135 0 0.176433f
c_60 XROM/XI7/XI4/NET99 0 0.176433f
c_61 XROM/XI7/XI4/NET127 0 0.176433f
c_62 XROM/XI7/XI4/NET91 0 0.176433f
c_63 XROM/XI7/XI4/NET119 0 0.176433f
c_64 XROM/XI7/XI4/NET83 0 0.136314f
c_65 XROM/XI6/XI3/NET143 0 0.14368f
c_66 XROM/XI6/XI3/NET107 0 0.176433f
c_67 XROM/XI6/XI3/NET135 0 0.176433f
c_68 XROM/XI6/XI3/NET99 0 0.176433f
c_69 XROM/XI6/XI3/NET127 0 0.176433f
c_70 XROM/XI6/XI3/NET91 0 0.176433f
c_71 XROM/XI6/XI3/NET119 0 0.176433f
c_72 XROM/XI6/XI3/NET83 0 0.176433f
c_73 XROM/XI6/XI7/NET143 0 0.176433f
c_74 XROM/XI6/XI7/NET107 0 0.176433f
c_75 XROM/XI6/XI7/NET135 0 0.176433f
c_76 XROM/XI6/XI7/NET99 0 0.176433f
c_77 XROM/XI6/XI7/NET127 0 0.176433f
c_78 XROM/XI6/XI7/NET91 0 0.176433f
c_79 XROM/XI6/XI7/NET119 0 0.176433f
c_80 XROM/XI6/XI7/NET83 0 0.136314f
c_81 XROM/XI6/XI2/NET143 0 0.138821f
c_82 XROM/XI6/XI2/NET107 0 0.176433f
c_83 XROM/XI6/XI2/NET135 0 0.176433f
c_84 XROM/XI6/XI2/NET99 0 0.176433f
c_85 XROM/XI6/XI2/NET127 0 0.176433f
c_86 XROM/XI6/XI2/NET91 0 0.176433f
c_87 XROM/XI6/XI2/NET119 0 0.176433f
c_88 XROM/XI6/XI2/NET83 0 0.176433f
c_89 XROM/XI6/XI6/NET143 0 0.176433f
c_90 XROM/XI6/XI6/NET107 0 0.176433f
c_91 XROM/XI6/XI6/NET135 0 0.176433f
c_92 XROM/XI6/XI6/NET99 0 0.176433f
c_93 XROM/XI6/XI6/NET127 0 0.176433f
c_94 XROM/XI6/XI6/NET91 0 0.176433f
c_95 XROM/XI6/XI6/NET119 0 0.176433f
c_96 XROM/XI6/XI6/NET83 0 0.136314f
c_97 XROM/XI6/XI1/NET143 0 0.142339f
c_98 XROM/XI6/XI1/NET107 0 0.176433f
c_99 XROM/XI6/XI1/NET135 0 0.176433f
c_100 XROM/XI6/XI1/NET99 0 0.176433f
c_101 XROM/XI6/XI1/NET127 0 0.176433f
c_102 XROM/XI6/XI1/NET91 0 0.176433f
c_103 XROM/XI6/XI1/NET119 0 0.176433f
c_104 XROM/XI6/XI1/NET83 0 0.176433f
c_105 XROM/XI6/XI5/NET143 0 0.176433f
c_106 XROM/XI6/XI5/NET107 0 0.176433f
c_107 XROM/XI6/XI5/NET135 0 0.176433f
c_108 XROM/XI6/XI5/NET99 0 0.176433f
c_109 XROM/XI6/XI5/NET127 0 0.176433f
c_110 XROM/XI6/XI5/NET91 0 0.176433f
c_111 XROM/XI6/XI5/NET119 0 0.176433f
c_112 XROM/XI6/XI5/NET83 0 0.136314f
c_113 XROM/XI6/XI0/NET143 0 0.14368f
c_114 XROM/XI6/XI0/NET107 0 0.176433f
c_115 XROM/XI6/XI0/NET135 0 0.176433f
c_116 XROM/XI6/XI0/NET99 0 0.176433f
c_117 XROM/XI6/XI0/NET127 0 0.176433f
c_118 XROM/XI6/XI0/NET91 0 0.176433f
c_119 XROM/XI6/XI0/NET119 0 0.176433f
c_120 XROM/XI6/XI0/NET83 0 0.176433f
c_121 XROM/XI6/XI4/NET143 0 0.176433f
c_122 XROM/XI6/XI4/NET107 0 0.176433f
c_123 XROM/XI6/XI4/NET135 0 0.176433f
c_124 XROM/XI6/XI4/NET99 0 0.176433f
c_125 XROM/XI6/XI4/NET127 0 0.176433f
c_126 XROM/XI6/XI4/NET91 0 0.176433f
c_127 XROM/XI6/XI4/NET119 0 0.176433f
c_128 XROM/XI6/XI4/NET83 0 0.136314f
c_129 XROM/XI5/XI3/NET143 0 0.14368f
c_130 XROM/XI5/XI3/NET107 0 0.18066f
c_131 XROM/XI5/XI3/NET135 0 0.176433f
c_132 XROM/XI5/XI3/NET99 0 0.18066f
c_133 XROM/XI5/XI3/NET127 0 0.176433f
c_134 XROM/XI5/XI3/NET91 0 0.18066f
c_135 XROM/XI5/XI3/NET119 0 0.176433f
c_136 XROM/XI5/XI3/NET83 0 0.18066f
c_137 XROM/XI5/XI7/NET143 0 0.176433f
c_138 XROM/XI5/XI7/NET107 0 0.18066f
c_139 XROM/XI5/XI7/NET135 0 0.176433f
c_140 XROM/XI5/XI7/NET99 0 0.18066f
c_141 XROM/XI5/XI7/NET127 0 0.176433f
c_142 XROM/XI5/XI7/NET91 0 0.18066f
c_143 XROM/XI5/XI7/NET119 0 0.176433f
c_144 XROM/XI5/XI7/NET83 0 0.138908f
c_145 XROM/XI5/XI2/NET143 0 0.138821f
c_146 XROM/XI5/XI2/NET107 0 0.176433f
c_147 XROM/XI5/XI2/NET135 0 0.176433f
c_148 XROM/XI5/XI2/NET99 0 0.176433f
c_149 XROM/XI5/XI2/NET127 0 0.176433f
c_150 XROM/XI5/XI2/NET91 0 0.176433f
c_151 XROM/XI5/XI2/NET119 0 0.176433f
c_152 XROM/XI5/XI2/NET83 0 0.176433f
c_153 XROM/XI5/XI6/NET143 0 0.176433f
c_154 XROM/XI5/XI6/NET107 0 0.176433f
c_155 XROM/XI5/XI6/NET135 0 0.176433f
c_156 XROM/XI5/XI6/NET99 0 0.176433f
c_157 XROM/XI5/XI6/NET127 0 0.176433f
c_158 XROM/XI5/XI6/NET91 0 0.176433f
c_159 XROM/XI5/XI6/NET119 0 0.176433f
c_160 XROM/XI5/XI6/NET83 0 0.136314f
c_161 XROM/XI5/XI1/NET143 0 0.142339f
c_162 XROM/XI5/XI1/NET107 0 0.176433f
c_163 XROM/XI5/XI1/NET135 0 0.176433f
c_164 XROM/XI5/XI1/NET99 0 0.176433f
c_165 XROM/XI5/XI1/NET127 0 0.176433f
c_166 XROM/XI5/XI1/NET91 0 0.176433f
c_167 XROM/XI5/XI1/NET119 0 0.176433f
c_168 XROM/XI5/XI1/NET83 0 0.176433f
c_169 XROM/XI5/XI5/NET143 0 0.176433f
c_170 XROM/XI5/XI5/NET107 0 0.176433f
c_171 XROM/XI5/XI5/NET135 0 0.176433f
c_172 XROM/XI5/XI5/NET99 0 0.176433f
c_173 XROM/XI5/XI5/NET127 0 0.176433f
c_174 XROM/XI5/XI5/NET91 0 0.176433f
c_175 XROM/XI5/XI5/NET119 0 0.176433f
c_176 XROM/XI5/XI5/NET83 0 0.136314f
c_177 XROM/XI5/XI0/NET143 0 0.14368f
c_178 XROM/XI5/XI0/NET107 0 0.176433f
c_179 XROM/XI5/XI0/NET135 0 0.176433f
c_180 XROM/XI5/XI0/NET99 0 0.176433f
c_181 XROM/XI5/XI0/NET127 0 0.176433f
c_182 XROM/XI5/XI0/NET91 0 0.176433f
c_183 XROM/XI5/XI0/NET119 0 0.176433f
c_184 XROM/XI5/XI0/NET83 0 0.176433f
c_185 XROM/XI5/XI4/NET143 0 0.176433f
c_186 XROM/XI5/XI4/NET107 0 0.176433f
c_187 XROM/XI5/XI4/NET135 0 0.176433f
c_188 XROM/XI5/XI4/NET99 0 0.176433f
c_189 XROM/XI5/XI4/NET127 0 0.176433f
c_190 XROM/XI5/XI4/NET91 0 0.176433f
c_191 XROM/XI5/XI4/NET119 0 0.176433f
c_192 XROM/XI5/XI4/NET83 0 0.136314f
c_193 XROM/XI4/XI3/NET143 0 0.14368f
c_194 XROM/XI4/XI3/NET107 0 0.176433f
c_195 XROM/XI4/XI3/NET135 0 0.176433f
c_196 XROM/XI4/XI3/NET99 0 0.176433f
c_197 XROM/XI4/XI3/NET127 0 0.176433f
c_198 XROM/XI4/XI3/NET91 0 0.176433f
c_199 XROM/XI4/XI3/NET119 0 0.176433f
c_200 XROM/XI4/XI3/NET83 0 0.176433f
c_201 XROM/XI4/XI7/NET143 0 0.176433f
c_202 XROM/XI4/XI7/NET107 0 0.176433f
c_203 XROM/XI4/XI7/NET135 0 0.176433f
c_204 XROM/XI4/XI7/NET99 0 0.176433f
c_205 XROM/XI4/XI7/NET127 0 0.176433f
c_206 XROM/XI4/XI7/NET91 0 0.176433f
c_207 XROM/XI4/XI7/NET119 0 0.176433f
c_208 XROM/XI4/XI7/NET83 0 0.136314f
c_209 XROM/XI4/XI2/NET143 0 0.138821f
c_210 XROM/XI4/XI2/NET107 0 0.176433f
c_211 XROM/XI4/XI2/NET135 0 0.176433f
c_212 XROM/XI4/XI2/NET99 0 0.176433f
c_213 XROM/XI4/XI2/NET127 0 0.176433f
c_214 XROM/XI4/XI2/NET91 0 0.176433f
c_215 XROM/XI4/XI2/NET119 0 0.176433f
c_216 XROM/XI4/XI2/NET83 0 0.176433f
c_217 XROM/XI4/XI6/NET143 0 0.176433f
c_218 XROM/XI4/XI6/NET107 0 0.176433f
c_219 XROM/XI4/XI6/NET135 0 0.176433f
c_220 XROM/XI4/XI6/NET99 0 0.176433f
c_221 XROM/XI4/XI6/NET127 0 0.176433f
c_222 XROM/XI4/XI6/NET91 0 0.176433f
c_223 XROM/XI4/XI6/NET119 0 0.176433f
c_224 XROM/XI4/XI6/NET83 0 0.136314f
c_225 XROM/XI4/XI1/NET143 0 0.142339f
c_226 XROM/XI4/XI1/NET107 0 0.176433f
c_227 XROM/XI4/XI1/NET135 0 0.176433f
c_228 XROM/XI4/XI1/NET99 0 0.176433f
c_229 XROM/XI4/XI1/NET127 0 0.176433f
c_230 XROM/XI4/XI1/NET91 0 0.176433f
c_231 XROM/XI4/XI1/NET119 0 0.176433f
c_232 XROM/XI4/XI1/NET83 0 0.176433f
c_233 XROM/XI4/XI5/NET143 0 0.176433f
c_234 XROM/XI4/XI5/NET107 0 0.176433f
c_235 XROM/XI4/XI5/NET135 0 0.176433f
c_236 XROM/XI4/XI5/NET99 0 0.176433f
c_237 XROM/XI4/XI5/NET127 0 0.176433f
c_238 XROM/XI4/XI5/NET91 0 0.176433f
c_239 XROM/XI4/XI5/NET119 0 0.176433f
c_240 XROM/XI4/XI5/NET83 0 0.136314f
c_241 XROM/XI4/XI0/NET143 0 0.14368f
c_242 XROM/XI4/XI0/NET107 0 0.176433f
c_243 XROM/XI4/XI0/NET135 0 0.176433f
c_244 XROM/XI4/XI0/NET99 0 0.176433f
c_245 XROM/XI4/XI0/NET127 0 0.176433f
c_246 XROM/XI4/XI0/NET91 0 0.176433f
c_247 XROM/XI4/XI0/NET119 0 0.176433f
c_248 XROM/XI4/XI0/NET83 0 0.176433f
c_249 XROM/XI4/XI4/NET143 0 0.176433f
c_250 XROM/XI4/XI4/NET107 0 0.176433f
c_251 XROM/XI4/XI4/NET135 0 0.176433f
c_252 XROM/XI4/XI4/NET99 0 0.176433f
c_253 XROM/XI4/XI4/NET127 0 0.176433f
c_254 XROM/XI4/XI4/NET91 0 0.176433f
c_255 XROM/XI4/XI4/NET119 0 0.176433f
c_256 XROM/XI4/XI4/NET83 0 0.136314f
c_257 XROM/XI3/XI3/NET143 0 0.14368f
c_258 XROM/XI3/XI3/NET107 0 0.18066f
c_259 XROM/XI3/XI3/NET135 0 0.176433f
c_260 XROM/XI3/XI3/NET99 0 0.18066f
c_261 XROM/XI3/XI3/NET127 0 0.176433f
c_262 XROM/XI3/XI3/NET91 0 0.18066f
c_263 XROM/XI3/XI3/NET119 0 0.176433f
c_264 XROM/XI3/XI3/NET83 0 0.18066f
c_265 XROM/XI3/XI7/NET143 0 0.176433f
c_266 XROM/XI3/XI7/NET107 0 0.18066f
c_267 XROM/XI3/XI7/NET135 0 0.176433f
c_268 XROM/XI3/XI7/NET99 0 0.18066f
c_269 XROM/XI3/XI7/NET127 0 0.176433f
c_270 XROM/XI3/XI7/NET91 0 0.18066f
c_271 XROM/XI3/XI7/NET119 0 0.176433f
c_272 XROM/XI3/XI7/NET83 0 0.138908f
c_273 XROM/XI3/XI2/NET143 0 0.138821f
c_274 XROM/XI3/XI2/NET107 0 0.176433f
c_275 XROM/XI3/XI2/NET135 0 0.176433f
c_276 XROM/XI3/XI2/NET99 0 0.176433f
c_277 XROM/XI3/XI2/NET127 0 0.176433f
c_278 XROM/XI3/XI2/NET91 0 0.176433f
c_279 XROM/XI3/XI2/NET119 0 0.176433f
c_280 XROM/XI3/XI2/NET83 0 0.176433f
c_281 XROM/XI3/XI6/NET143 0 0.176433f
c_282 XROM/XI3/XI6/NET107 0 0.176433f
c_283 XROM/XI3/XI6/NET135 0 0.176433f
c_284 XROM/XI3/XI6/NET99 0 0.176433f
c_285 XROM/XI3/XI6/NET127 0 0.176433f
c_286 XROM/XI3/XI6/NET91 0 0.176433f
c_287 XROM/XI3/XI6/NET119 0 0.176433f
c_288 XROM/XI3/XI6/NET83 0 0.136314f
c_289 XROM/XI3/XI1/NET143 0 0.142339f
c_290 XROM/XI3/XI1/NET107 0 0.176433f
c_291 XROM/XI3/XI1/NET135 0 0.176433f
c_292 XROM/XI3/XI1/NET99 0 0.176433f
c_293 XROM/XI3/XI1/NET127 0 0.176433f
c_294 XROM/XI3/XI1/NET91 0 0.176433f
c_295 XROM/XI3/XI1/NET119 0 0.176433f
c_296 XROM/XI3/XI1/NET83 0 0.176433f
c_297 XROM/XI3/XI5/NET143 0 0.176433f
c_298 XROM/XI3/XI5/NET107 0 0.176433f
c_299 XROM/XI3/XI5/NET135 0 0.176433f
c_300 XROM/XI3/XI5/NET99 0 0.176433f
c_301 XROM/XI3/XI5/NET127 0 0.176433f
c_302 XROM/XI3/XI5/NET91 0 0.176433f
c_303 XROM/XI3/XI5/NET119 0 0.176433f
c_304 XROM/XI3/XI5/NET83 0 0.136314f
c_305 XROM/XI3/XI0/NET143 0 0.14368f
c_306 XROM/XI3/XI0/NET107 0 0.176433f
c_307 XROM/XI3/XI0/NET135 0 0.176433f
c_308 XROM/XI3/XI0/NET99 0 0.176433f
c_309 XROM/XI3/XI0/NET127 0 0.176433f
c_310 XROM/XI3/XI0/NET91 0 0.176433f
c_311 XROM/XI3/XI0/NET119 0 0.176433f
c_312 XROM/XI3/XI0/NET83 0 0.176433f
c_313 XROM/XI3/XI4/NET143 0 0.176433f
c_314 XROM/XI3/XI4/NET107 0 0.176433f
c_315 XROM/XI3/XI4/NET135 0 0.176433f
c_316 XROM/XI3/XI4/NET99 0 0.176433f
c_317 XROM/XI3/XI4/NET127 0 0.176433f
c_318 XROM/XI3/XI4/NET91 0 0.176433f
c_319 XROM/XI3/XI4/NET119 0 0.176433f
c_320 XROM/XI3/XI4/NET83 0 0.136314f
c_321 XROM/XI2/XI3/NET143 0 0.14368f
c_322 XROM/XI2/XI3/NET107 0 0.176433f
c_323 XROM/XI2/XI3/NET135 0 0.176433f
c_324 XROM/XI2/XI3/NET99 0 0.176433f
c_325 XROM/XI2/XI3/NET127 0 0.176433f
c_326 XROM/XI2/XI3/NET91 0 0.176433f
c_327 XROM/XI2/XI3/NET119 0 0.176433f
c_328 XROM/XI2/XI3/NET83 0 0.176433f
c_329 XROM/XI2/XI7/NET143 0 0.176433f
c_330 XROM/XI2/XI7/NET107 0 0.176433f
c_331 XROM/XI2/XI7/NET135 0 0.176433f
c_332 XROM/XI2/XI7/NET99 0 0.176433f
c_333 XROM/XI2/XI7/NET127 0 0.176433f
c_334 XROM/XI2/XI7/NET91 0 0.176433f
c_335 XROM/XI2/XI7/NET119 0 0.176433f
c_336 XROM/XI2/XI7/NET83 0 0.136314f
c_337 XROM/XI2/XI2/NET143 0 0.138821f
c_338 XROM/XI2/XI2/NET107 0 0.176433f
c_339 XROM/XI2/XI2/NET135 0 0.176433f
c_340 XROM/XI2/XI2/NET99 0 0.176433f
c_341 XROM/XI2/XI2/NET127 0 0.176433f
c_342 XROM/XI2/XI2/NET91 0 0.176433f
c_343 XROM/XI2/XI2/NET119 0 0.176433f
c_344 XROM/XI2/XI2/NET83 0 0.176433f
c_345 XROM/XI2/XI6/NET143 0 0.176433f
c_346 XROM/XI2/XI6/NET107 0 0.176433f
c_347 XROM/XI2/XI6/NET135 0 0.176433f
c_348 XROM/XI2/XI6/NET99 0 0.176433f
c_349 XROM/XI2/XI6/NET127 0 0.176433f
c_350 XROM/XI2/XI6/NET91 0 0.176433f
c_351 XROM/XI2/XI6/NET119 0 0.176433f
c_352 XROM/XI2/XI6/NET83 0 0.136314f
c_353 XROM/XI2/XI1/NET143 0 0.142339f
c_354 XROM/XI2/XI1/NET107 0 0.176433f
c_355 XROM/XI2/XI1/NET135 0 0.176433f
c_356 XROM/XI2/XI1/NET99 0 0.176433f
c_357 XROM/XI2/XI1/NET127 0 0.176433f
c_358 XROM/XI2/XI1/NET91 0 0.176433f
c_359 XROM/XI2/XI1/NET119 0 0.176433f
c_360 XROM/XI2/XI1/NET83 0 0.176433f
c_361 XROM/XI2/XI5/NET143 0 0.176433f
c_362 XROM/XI2/XI5/NET107 0 0.176433f
c_363 XROM/XI2/XI5/NET135 0 0.176433f
c_364 XROM/XI2/XI5/NET99 0 0.176433f
c_365 XROM/XI2/XI5/NET127 0 0.176433f
c_366 XROM/XI2/XI5/NET91 0 0.176433f
c_367 XROM/XI2/XI5/NET119 0 0.176433f
c_368 XROM/XI2/XI5/NET83 0 0.136314f
c_369 XROM/XI2/XI0/NET143 0 0.14368f
c_370 XROM/XI2/XI0/NET107 0 0.176433f
c_371 XROM/XI2/XI0/NET135 0 0.176433f
c_372 XROM/XI2/XI0/NET99 0 0.176433f
c_373 XROM/XI2/XI0/NET127 0 0.176433f
c_374 XROM/XI2/XI0/NET91 0 0.176433f
c_375 XROM/XI2/XI0/NET119 0 0.176433f
c_376 XROM/XI2/XI0/NET83 0 0.176433f
c_377 XROM/XI2/XI4/NET143 0 0.176433f
c_378 XROM/XI2/XI4/NET107 0 0.176433f
c_379 XROM/XI2/XI4/NET135 0 0.176433f
c_380 XROM/XI2/XI4/NET99 0 0.176433f
c_381 XROM/XI2/XI4/NET127 0 0.176433f
c_382 XROM/XI2/XI4/NET91 0 0.176433f
c_383 XROM/XI2/XI4/NET119 0 0.176433f
c_384 XROM/XI2/XI4/NET83 0 0.136314f
c_385 XROM/XI1/XI3/NET143 0 0.14368f
c_386 XROM/XI1/XI3/NET107 0 0.18066f
c_387 XROM/XI1/XI3/NET135 0 0.176433f
c_388 XROM/XI1/XI3/NET99 0 0.18066f
c_389 XROM/XI1/XI3/NET127 0 0.176433f
c_390 XROM/XI1/XI3/NET91 0 0.18066f
c_391 XROM/XI1/XI3/NET119 0 0.176433f
c_392 XROM/XI1/XI3/NET83 0 0.18066f
c_393 XROM/XI1/XI7/NET143 0 0.176433f
c_394 XROM/XI1/XI7/NET107 0 0.18066f
c_395 XROM/XI1/XI7/NET135 0 0.176433f
c_396 XROM/XI1/XI7/NET99 0 0.18066f
c_397 XROM/XI1/XI7/NET127 0 0.176433f
c_398 XROM/XI1/XI7/NET83 0 0.18066f
c_399 XROM/XI1/XI7/NET119 0 0.176433f
c_400 XROM/XI1/XI7/NET91 0 0.138908f
c_401 XROM/XI1/XI2/NET143 0 0.138821f
c_402 XROM/XI1/XI2/NET107 0 0.176433f
c_403 XROM/XI1/XI2/NET135 0 0.176433f
c_404 XROM/XI1/XI2/NET99 0 0.176433f
c_405 XROM/XI1/XI2/NET127 0 0.176433f
c_406 XROM/XI1/XI2/NET91 0 0.176433f
c_407 XROM/XI1/XI2/NET119 0 0.176433f
c_408 XROM/XI1/XI2/NET83 0 0.176433f
c_409 XROM/XI1/XI6/NET143 0 0.176433f
c_410 XROM/XI1/XI6/NET107 0 0.176433f
c_411 XROM/XI1/XI6/NET135 0 0.176433f
c_412 XROM/XI1/XI6/NET99 0 0.176433f
c_413 XROM/XI1/XI6/NET127 0 0.176433f
c_414 XROM/XI1/XI6/NET83 0 0.176433f
c_415 XROM/XI1/XI6/NET119 0 0.176433f
c_416 XROM/XI1/XI6/NET91 0 0.136314f
c_417 XROM/XI1/XI1/NET143 0 0.142339f
c_418 XROM/XI1/XI1/NET107 0 0.176433f
c_419 XROM/XI1/XI1/NET135 0 0.176433f
c_420 XROM/XI1/XI1/NET99 0 0.176433f
c_421 XROM/XI1/XI1/NET127 0 0.176433f
c_422 XROM/XI1/XI1/NET91 0 0.176433f
c_423 XROM/XI1/XI1/NET119 0 0.176433f
c_424 XROM/XI1/XI1/NET83 0 0.176433f
c_425 XROM/XI1/XI5/NET143 0 0.176433f
c_426 XROM/XI1/XI5/NET107 0 0.176433f
c_427 XROM/XI1/XI5/NET135 0 0.176433f
c_428 XROM/XI1/XI5/NET99 0 0.176433f
c_429 XROM/XI1/XI5/NET127 0 0.176433f
c_430 XROM/XI1/XI5/NET83 0 0.176433f
c_431 XROM/XI1/XI5/NET119 0 0.176433f
c_432 XROM/XI1/XI5/NET91 0 0.136314f
c_433 XROM/XI1/XI0/NET143 0 0.14368f
c_434 XROM/XI1/XI0/NET107 0 0.176433f
c_435 XROM/XI1/XI0/NET135 0 0.176433f
c_436 XROM/XI1/XI0/NET99 0 0.176433f
c_437 XROM/XI1/XI0/NET127 0 0.176433f
c_438 XROM/XI1/XI0/NET91 0 0.176433f
c_439 XROM/XI1/XI0/NET119 0 0.176433f
c_440 XROM/XI1/XI0/NET83 0 0.176433f
c_441 XROM/XI1/XI4/NET143 0 0.176433f
c_442 XROM/XI1/XI4/NET107 0 0.176433f
c_443 XROM/XI1/XI4/NET135 0 0.176433f
c_444 XROM/XI1/XI4/NET99 0 0.176433f
c_445 XROM/XI1/XI4/NET127 0 0.176433f
c_446 XROM/XI1/XI4/NET83 0 0.176433f
c_447 XROM/XI1/XI4/NET119 0 0.176433f
c_448 XROM/XI1/XI4/NET91 0 0.136314f
c_449 XROM/XI0/XI3/NET143 0 0.14368f
c_450 XROM/XI0/XI3/NET107 0 0.176433f
c_451 XROM/XI0/XI3/NET135 0 0.176433f
c_452 XROM/XI0/XI3/NET99 0 0.176433f
c_453 XROM/XI0/XI3/NET127 0 0.176433f
c_454 XROM/XI0/XI3/NET91 0 0.176433f
c_455 XROM/XI0/XI3/NET119 0 0.176433f
c_456 XROM/XI0/XI3/NET83 0 0.176433f
c_457 XROM/XI0/XI7/NET143 0 0.176433f
c_458 XROM/XI0/XI7/NET107 0 0.176433f
c_459 XROM/XI0/XI7/NET135 0 0.176433f
c_460 XROM/XI0/XI7/NET99 0 0.176433f
c_461 XROM/XI0/XI7/NET127 0 0.176433f
c_462 XROM/XI0/XI7/NET83 0 0.176433f
c_463 XROM/XI0/XI7/NET119 0 0.176433f
c_464 XROM/XI0/XI7/NET91 0 0.136314f
c_465 XROM/XI0/XI2/NET143 0 0.138821f
c_466 XROM/XI0/XI2/NET107 0 0.176433f
c_467 XROM/XI0/XI2/NET135 0 0.176433f
c_468 XROM/XI0/XI2/NET99 0 0.176433f
c_469 XROM/XI0/XI2/NET127 0 0.176433f
c_470 XROM/XI0/XI2/NET91 0 0.176433f
c_471 XROM/XI0/XI2/NET119 0 0.176433f
c_472 XROM/XI0/XI2/NET83 0 0.176433f
c_473 XROM/XI0/XI6/NET143 0 0.176433f
c_474 XROM/XI0/XI6/NET107 0 0.176433f
c_475 XROM/XI0/XI6/NET135 0 0.176433f
c_476 XROM/XI0/XI6/NET91 0 0.176433f
c_477 XROM/XI0/XI6/NET119 0 0.176433f
c_478 XROM/XI0/XI6/NET83 0 0.176433f
c_479 XROM/XI0/XI6/NET127 0 0.176433f
c_480 XROM/XI0/XI6/NET99 0 0.136314f
c_481 XROM/XI0/XI1/NET143 0 0.142339f
c_482 XROM/XI0/XI1/NET107 0 0.176433f
c_483 XROM/XI0/XI1/NET135 0 0.176433f
c_484 XROM/XI0/XI1/NET99 0 0.176433f
c_485 XROM/XI0/XI1/NET127 0 0.176433f
c_486 XROM/XI0/XI1/NET91 0 0.176433f
c_487 XROM/XI0/XI1/NET119 0 0.176433f
c_488 XROM/XI0/XI1/NET83 0 0.176433f
c_489 XROM/XI0/XI5/NET143 0 0.176433f
c_490 XROM/XI0/XI5/NET107 0 0.176433f
c_491 XROM/XI0/XI5/NET135 0 0.176433f
c_492 XROM/XI0/XI5/NET91 0 0.176433f
c_493 XROM/XI0/XI5/NET119 0 0.176433f
c_494 XROM/XI0/XI5/NET83 0 0.176433f
c_495 XROM/XI0/XI5/NET127 0 0.176433f
c_496 XROM/XI0/XI5/NET99 0 0.136314f
c_497 XROM/XI0/XI0/NET143 0 0.14368f
c_498 XROM/XI0/XI0/NET107 0 0.176433f
c_499 XROM/XI0/XI0/NET135 0 0.176433f
c_500 XROM/XI0/XI0/NET99 0 0.176433f
c_501 XROM/XI0/XI0/NET127 0 0.176433f
c_502 XROM/XI0/XI0/NET91 0 0.176433f
c_503 XROM/XI0/XI0/NET119 0 0.176433f
c_504 XROM/XI0/XI0/NET83 0 0.176433f
c_505 XROM/XI0/XI4/NET143 0 0.176433f
c_506 XROM/XI0/XI4/NET107 0 0.176433f
c_507 XROM/XI0/XI4/NET135 0 0.176433f
c_508 XROM/XI0/XI4/NET91 0 0.176433f
c_509 XROM/XI0/XI4/NET119 0 0.176433f
c_510 XROM/XI0/XI4/NET83 0 0.176433f
c_511 XROM/XI0/XI4/NET127 0 0.176433f
c_512 XROM/XI0/XI4/NET99 0 0.136314f
*
.include "top.pex.spi.TOP.pxi"
*
.ends
*
*
