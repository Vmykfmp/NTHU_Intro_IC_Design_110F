* SPICE NETLIST
***************************************
*HW2_Inverter_Chain_Branch_postsim
.lib 'cic018.l' TT
.temp 25
.unprot
.inc "ICB.pex.spi"
.option post

*Voltage
V1 VDD 0 1.8
V2 GND 0 0
VVIN_pulse VIN gnd pulse 0 1.8 10n 1n 1n 4n 10n

*Capacitor
CLa Vaout gnd 10pF
CLb Vbout gnd 10pF
CLc Vcout gnd 10pF

*Circuit
x1 GND VDD Vin Vaout Vbout Vcout ICB

*simulation setup
.Tran 1ps 50ns
.MEAS tran TpHL_N2 trig V(Vin) val=0.9 td=0 rise=1 targ V(Vaout) val=0.9 fall=1
.MEAS tran TpLH_N2 trig V(Vin) val=0.9 td=0 fall=1 targ V(Vaout) val=0.9 rise=1

.MEAS tran TpHL_N4 trig V(Vin) val=0.9 td=0 rise=1 targ V(Vbout) val=0.9 fall=1
.MEAS tran TpLH_N4 trig V(Vin) val=0.9 td=0 fall=1 targ V(Vbout) val=0.9 rise=1

.MEAS tran TpLL_N8 trig V(Vin) val=0.9 td=0 rise=1 targ V(Vcout) val=0.9 fall=1
.MEAS tran TpHH_N8 trig V(Vin) val=0.9 td=0 fall=1 targ V(Vcout) val=0.9 rise=1

.SUBCKT L POS NEG
.ENDS
.end
***************************************
.SUBCKT ICB GND VDD Vin Vaout Vbout Vcout
** N=20 EP=6 IP=0 FDC=3566
M0 4 Vin GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=-145 $Y=-166 $D=0
M1 5 4 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=1415 $Y=-166 $D=0
M2 GND 4 5 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=2105 $Y=-166 $D=0
M3 5 4 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=2795 $Y=-166 $D=0
M4 GND 4 5 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=3485 $Y=-166 $D=0
M5 5 4 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=4175 $Y=-166 $D=0
M6 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=5735 $Y=-166 $D=0
M7 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=6425 $Y=-166 $D=0
M8 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=7115 $Y=-166 $D=0
M9 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=7805 $Y=-166 $D=0
M10 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=8495 $Y=-166 $D=0
M11 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=9185 $Y=-166 $D=0
M12 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=9875 $Y=-166 $D=0
M13 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=10565 $Y=-166 $D=0
M14 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=11255 $Y=-166 $D=0
M15 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=11945 $Y=-166 $D=0
M16 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=12635 $Y=-166 $D=0
M17 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=13325 $Y=-166 $D=0
M18 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=14015 $Y=-166 $D=0
M19 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=14705 $Y=-166 $D=0
M20 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=15395 $Y=-166 $D=0
M21 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=16085 $Y=-166 $D=0
M22 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=16775 $Y=-166 $D=0
M23 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=17465 $Y=-166 $D=0
M24 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=18155 $Y=-166 $D=0
M25 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=18845 $Y=-166 $D=0
M26 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=19535 $Y=-166 $D=0
M27 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=20225 $Y=-166 $D=0
M28 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=20915 $Y=-166 $D=0
M29 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=21605 $Y=-166 $D=0
M30 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=22295 $Y=-166 $D=0
M31 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=22985 $Y=-166 $D=0
M32 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=23675 $Y=-166 $D=0
M33 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=24365 $Y=-166 $D=0
M34 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=25055 $Y=-166 $D=0
M35 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=25745 $Y=-166 $D=0
M36 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=26435 $Y=-166 $D=0
M37 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=27125 $Y=-166 $D=0
M38 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=27815 $Y=-166 $D=0
M39 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=28505 $Y=-166 $D=0
M40 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=29195 $Y=-166 $D=0
M41 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=29885 $Y=-166 $D=0
M42 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=30575 $Y=-166 $D=0
M43 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=31265 $Y=-166 $D=0
M44 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=31955 $Y=-166 $D=0
M45 GND 5 6 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=32645 $Y=-166 $D=0
M46 6 5 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=33335 $Y=-166 $D=0
M47 7 6 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=38665 $Y=-7792 $D=0
M48 8 6 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=38665 $Y=-166 $D=0
M49 9 6 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06 $X=38665 $Y=7460 $D=0
M50 10 7 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=40225 $Y=-7792 $D=0
M51 11 8 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=40225 $Y=-166 $D=0
M52 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=40225 $Y=7460 $D=0
M53 GND 7 10 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=40915 $Y=-7792 $D=0
M54 GND 8 11 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=40915 $Y=-166 $D=0
M55 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=40915 $Y=7460 $D=0
M56 10 7 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=41605 $Y=-7792 $D=0
M57 11 8 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=41605 $Y=-166 $D=0
M58 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=41605 $Y=7460 $D=0
M59 GND 8 11 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=42295 $Y=-166 $D=0
M60 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=42295 $Y=7460 $D=0
M61 11 8 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=42985 $Y=-166 $D=0
M62 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=42985 $Y=7460 $D=0
M63 12 10 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=43165 $Y=-7792 $D=0
M64 GND 8 11 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=43675 $Y=-166 $D=0
M65 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=43675 $Y=7460 $D=0
M66 GND 10 12 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=43855 $Y=-7792 $D=0
M67 11 8 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=44365 $Y=-166 $D=0
M68 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=44365 $Y=7460 $D=0
M69 12 10 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=44545 $Y=-7792 $D=0
M70 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=45055 $Y=7460 $D=0
M71 GND 10 12 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=45235 $Y=-7792 $D=0
M72 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=45745 $Y=7460 $D=0
M73 12 10 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=45925 $Y=-7792 $D=0
M74 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=45925 $Y=-166 $D=0
M75 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=46435 $Y=7460 $D=0
M76 GND 10 12 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=46615 $Y=-7792 $D=0
M77 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=46615 $Y=-166 $D=0
M78 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=47125 $Y=7460 $D=0
M79 12 10 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=47305 $Y=-7792 $D=0
M80 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=47305 $Y=-166 $D=0
M81 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=47815 $Y=7460 $D=0
M82 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=47995 $Y=-166 $D=0
M83 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=48505 $Y=7460 $D=0
M84 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=48685 $Y=-166 $D=0
M85 13 12 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=48865 $Y=-7792 $D=0
M86 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=49195 $Y=7460 $D=0
M87 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=49375 $Y=-166 $D=0
M88 GND 12 13 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=49555 $Y=-7792 $D=0
M89 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=49885 $Y=7460 $D=0
M90 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=50065 $Y=-166 $D=0
M91 13 12 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=50245 $Y=-7792 $D=0
M92 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=50575 $Y=7460 $D=0
M93 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=50755 $Y=-166 $D=0
M94 GND 12 13 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=50935 $Y=-7792 $D=0
M95 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=51265 $Y=7460 $D=0
M96 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=51445 $Y=-166 $D=0
M97 13 12 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=51625 $Y=-7792 $D=0
M98 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=51955 $Y=7460 $D=0
M99 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=52135 $Y=-166 $D=0
M100 GND 12 13 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=52315 $Y=-7792 $D=0
M101 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=52645 $Y=7460 $D=0
M102 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=52825 $Y=-166 $D=0
M103 13 12 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=53005 $Y=-7792 $D=0
M104 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=53335 $Y=7460 $D=0
M105 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=53515 $Y=-166 $D=0
M106 GND 12 13 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=53695 $Y=-7792 $D=0
M107 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=54025 $Y=7460 $D=0
M108 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=54205 $Y=-166 $D=0
M109 13 12 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=54385 $Y=-7792 $D=0
M110 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=54715 $Y=7460 $D=0
M111 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=54895 $Y=-166 $D=0
M112 GND 12 13 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=55075 $Y=-7792 $D=0
M113 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=55405 $Y=7460 $D=0
M114 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=55585 $Y=-166 $D=0
M115 13 12 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=55765 $Y=-7792 $D=0
M116 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=56095 $Y=7460 $D=0
M117 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=56275 $Y=-166 $D=0
M118 GND 12 13 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=56455 $Y=-7792 $D=0
M119 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=56785 $Y=7460 $D=0
M120 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=56965 $Y=-166 $D=0
M121 13 12 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=57145 $Y=-7792 $D=0
M122 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=57475 $Y=7460 $D=0
M123 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=57655 $Y=-166 $D=0
M124 GND 12 13 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=57835 $Y=-7792 $D=0
M125 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=58165 $Y=7460 $D=0
M126 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=58345 $Y=-166 $D=0
M127 13 12 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=58525 $Y=-7792 $D=0
M128 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=58855 $Y=7460 $D=0
M129 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=59035 $Y=-166 $D=0
M130 GND 12 13 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=59215 $Y=-7792 $D=0
M131 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=59545 $Y=7460 $D=0
M132 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=59725 $Y=-166 $D=0
M133 13 12 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=59905 $Y=-7792 $D=0
M134 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=60235 $Y=7460 $D=0
M135 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=60415 $Y=-166 $D=0
M136 GND 12 13 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=60595 $Y=-7792 $D=0
M137 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=60925 $Y=7460 $D=0
M138 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=61105 $Y=-166 $D=0
M139 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=61615 $Y=7460 $D=0
M140 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=61795 $Y=-166 $D=0
M141 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=62155 $Y=-7792 $D=0
M142 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=62305 $Y=7460 $D=0
M143 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=62485 $Y=-166 $D=0
M144 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=62845 $Y=-7792 $D=0
M145 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=62995 $Y=7460 $D=0
M146 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=63175 $Y=-166 $D=0
M147 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=63535 $Y=-7792 $D=0
M148 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=63685 $Y=7460 $D=0
M149 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=63865 $Y=-166 $D=0
M150 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=64225 $Y=-7792 $D=0
M151 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=64375 $Y=7460 $D=0
M152 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=64555 $Y=-166 $D=0
M153 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=64915 $Y=-7792 $D=0
M154 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=65065 $Y=7460 $D=0
M155 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=65245 $Y=-166 $D=0
M156 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=65605 $Y=-7792 $D=0
M157 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=65755 $Y=7460 $D=0
M158 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=65935 $Y=-166 $D=0
M159 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=66295 $Y=-7792 $D=0
M160 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=66445 $Y=7460 $D=0
M161 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=66625 $Y=-166 $D=0
M162 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=66985 $Y=-7792 $D=0
M163 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=67135 $Y=7460 $D=0
M164 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=67315 $Y=-166 $D=0
M165 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=67675 $Y=-7792 $D=0
M166 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=67825 $Y=7460 $D=0
M167 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=68005 $Y=-166 $D=0
M168 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=68365 $Y=-7792 $D=0
M169 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=68515 $Y=7460 $D=0
M170 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=68695 $Y=-166 $D=0
M171 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=69055 $Y=-7792 $D=0
M172 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=69205 $Y=7460 $D=0
M173 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=69385 $Y=-166 $D=0
M174 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=69745 $Y=-7792 $D=0
M175 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=69895 $Y=7460 $D=0
M176 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=70075 $Y=-166 $D=0
M177 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=70435 $Y=-7792 $D=0
M178 Vaout 9 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=70585 $Y=7460 $D=0
M179 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=70765 $Y=-166 $D=0
M180 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=71125 $Y=-7792 $D=0
M181 GND 9 Vaout GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=71275 $Y=7460 $D=0
M182 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=71455 $Y=-166 $D=0
M183 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=71815 $Y=-7792 $D=0
M184 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=72145 $Y=-166 $D=0
M185 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=72505 $Y=-7792 $D=0
M186 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=72835 $Y=-166 $D=0
M187 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=73195 $Y=-7792 $D=0
M188 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=73525 $Y=-166 $D=0
M189 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=73885 $Y=-7792 $D=0
M190 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=74215 $Y=-166 $D=0
M191 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=74575 $Y=-7792 $D=0
M192 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=74905 $Y=-166 $D=0
M193 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=75265 $Y=-7792 $D=0
M194 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=75595 $Y=-166 $D=0
M195 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=75955 $Y=-7792 $D=0
M196 15 11 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=76285 $Y=-166 $D=0
M197 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=76645 $Y=-7792 $D=0
M198 GND 11 15 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=76975 $Y=-166 $D=0
M199 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=77335 $Y=-7792 $D=0
M200 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=78025 $Y=-7792 $D=0
M201 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=78535 $Y=-166 $D=0
M202 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=78715 $Y=-7792 $D=0
M203 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=79225 $Y=-166 $D=0
M204 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=79405 $Y=-7792 $D=0
M205 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=79915 $Y=-166 $D=0
M206 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=80095 $Y=-7792 $D=0
M207 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=80605 $Y=-166 $D=0
M208 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=80785 $Y=-7792 $D=0
M209 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=81295 $Y=-166 $D=0
M210 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=81475 $Y=-7792 $D=0
M211 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=81985 $Y=-166 $D=0
M212 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=82165 $Y=-7792 $D=0
M213 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=82675 $Y=-166 $D=0
M214 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=82855 $Y=-7792 $D=0
M215 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=83365 $Y=-166 $D=0
M216 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=83545 $Y=-7792 $D=0
M217 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=84055 $Y=-166 $D=0
M218 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=84235 $Y=-7792 $D=0
M219 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=84745 $Y=-166 $D=0
M220 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=84925 $Y=-7792 $D=0
M221 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=85435 $Y=-166 $D=0
M222 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=85615 $Y=-7792 $D=0
M223 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=86125 $Y=-166 $D=0
M224 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=86305 $Y=-7792 $D=0
M225 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=86815 $Y=-166 $D=0
M226 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=86995 $Y=-7792 $D=0
M227 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=87505 $Y=-166 $D=0
M228 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=87685 $Y=-7792 $D=0
M229 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=88195 $Y=-166 $D=0
M230 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=88375 $Y=-7792 $D=0
M231 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=88885 $Y=-166 $D=0
M232 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=89065 $Y=-7792 $D=0
M233 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=89575 $Y=-166 $D=0
M234 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=89755 $Y=-7792 $D=0
M235 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=90265 $Y=-166 $D=0
M236 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=90445 $Y=-7792 $D=0
M237 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=90955 $Y=-166 $D=0
M238 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=91135 $Y=-7792 $D=0
M239 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=91645 $Y=-166 $D=0
M240 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=91825 $Y=-7792 $D=0
M241 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=92335 $Y=-166 $D=0
M242 16 13 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=92515 $Y=-7792 $D=0
M243 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=93025 $Y=-166 $D=0
M244 GND 13 16 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=93205 $Y=-7792 $D=0
M245 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=93715 $Y=-166 $D=0
M246 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=94405 $Y=-166 $D=0
M247 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=94765 $Y=-7792 $D=0
M248 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=95095 $Y=-166 $D=0
M249 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=95455 $Y=-7792 $D=0
M250 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=95785 $Y=-166 $D=0
M251 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=96145 $Y=-7792 $D=0
M252 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=96475 $Y=-166 $D=0
M253 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=96835 $Y=-7792 $D=0
M254 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=97165 $Y=-166 $D=0
M255 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=97525 $Y=-7792 $D=0
M256 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=97855 $Y=-166 $D=0
M257 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=98215 $Y=-7792 $D=0
M258 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=98545 $Y=-166 $D=0
M259 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=98905 $Y=-7792 $D=0
M260 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=99235 $Y=-166 $D=0
M261 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=99595 $Y=-7792 $D=0
M262 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=99925 $Y=-166 $D=0
M263 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=100285 $Y=-7792 $D=0
M264 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=100615 $Y=-166 $D=0
M265 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=100975 $Y=-7792 $D=0
M266 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=101305 $Y=-166 $D=0
M267 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=101665 $Y=-7792 $D=0
M268 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=101995 $Y=-166 $D=0
M269 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=102355 $Y=-7792 $D=0
M270 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=102685 $Y=-166 $D=0
M271 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=103045 $Y=-7792 $D=0
M272 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=103375 $Y=-166 $D=0
M273 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=103735 $Y=-7792 $D=0
M274 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=104065 $Y=-166 $D=0
M275 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=104425 $Y=-7792 $D=0
M276 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=104755 $Y=-166 $D=0
M277 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=105115 $Y=-7792 $D=0
M278 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=105445 $Y=-166 $D=0
M279 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=105805 $Y=-7792 $D=0
M280 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=106135 $Y=-166 $D=0
M281 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=106495 $Y=-7792 $D=0
M282 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=106825 $Y=-166 $D=0
M283 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=107185 $Y=-7792 $D=0
M284 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=107515 $Y=-166 $D=0
M285 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=107875 $Y=-7792 $D=0
M286 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=108205 $Y=-166 $D=0
M287 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=108565 $Y=-7792 $D=0
M288 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=108895 $Y=-166 $D=0
M289 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=109255 $Y=-7792 $D=0
M290 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=109585 $Y=-166 $D=0
M291 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=109945 $Y=-7792 $D=0
M292 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=110275 $Y=-166 $D=0
M293 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=110635 $Y=-7792 $D=0
M294 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=110965 $Y=-166 $D=0
M295 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=111325 $Y=-7792 $D=0
M296 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=111655 $Y=-166 $D=0
M297 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=112015 $Y=-7792 $D=0
M298 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=112345 $Y=-166 $D=0
M299 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=112705 $Y=-7792 $D=0
M300 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=113035 $Y=-166 $D=0
M301 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=113395 $Y=-7792 $D=0
M302 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=113725 $Y=-166 $D=0
M303 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=114085 $Y=-7792 $D=0
M304 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=114415 $Y=-166 $D=0
M305 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=114775 $Y=-7792 $D=0
M306 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=115105 $Y=-166 $D=0
M307 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=115465 $Y=-7792 $D=0
M308 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=115795 $Y=-166 $D=0
M309 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=116155 $Y=-7792 $D=0
M310 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=116485 $Y=-166 $D=0
M311 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=116845 $Y=-7792 $D=0
M312 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=117175 $Y=-166 $D=0
M313 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=117535 $Y=-7792 $D=0
M314 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=117865 $Y=-166 $D=0
M315 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=118225 $Y=-7792 $D=0
M316 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=118555 $Y=-166 $D=0
M317 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=118915 $Y=-7792 $D=0
M318 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=119245 $Y=-166 $D=0
M319 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=119605 $Y=-7792 $D=0
M320 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=119935 $Y=-166 $D=0
M321 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=120295 $Y=-7792 $D=0
M322 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=120625 $Y=-166 $D=0
M323 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=120985 $Y=-7792 $D=0
M324 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=121315 $Y=-166 $D=0
M325 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=121675 $Y=-7792 $D=0
M326 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=122005 $Y=-166 $D=0
M327 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=122365 $Y=-7792 $D=0
M328 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=122695 $Y=-166 $D=0
M329 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=123055 $Y=-7792 $D=0
M330 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=123385 $Y=-166 $D=0
M331 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=123745 $Y=-7792 $D=0
M332 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=124075 $Y=-166 $D=0
M333 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=124435 $Y=-7792 $D=0
M334 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=124765 $Y=-166 $D=0
M335 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=125125 $Y=-7792 $D=0
M336 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=125455 $Y=-166 $D=0
M337 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=125815 $Y=-7792 $D=0
M338 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=126145 $Y=-166 $D=0
M339 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=126505 $Y=-7792 $D=0
M340 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=126835 $Y=-166 $D=0
M341 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=127195 $Y=-7792 $D=0
M342 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=127525 $Y=-166 $D=0
M343 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=127885 $Y=-7792 $D=0
M344 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=128215 $Y=-166 $D=0
M345 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=128575 $Y=-7792 $D=0
M346 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=128905 $Y=-166 $D=0
M347 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=129265 $Y=-7792 $D=0
M348 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=129595 $Y=-166 $D=0
M349 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=129955 $Y=-7792 $D=0
M350 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=130285 $Y=-166 $D=0
M351 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=130645 $Y=-7792 $D=0
M352 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=130975 $Y=-166 $D=0
M353 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=131335 $Y=-7792 $D=0
M354 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=131665 $Y=-166 $D=0
M355 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=132025 $Y=-7792 $D=0
M356 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=132355 $Y=-166 $D=0
M357 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=132715 $Y=-7792 $D=0
M358 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=133045 $Y=-166 $D=0
M359 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=133405 $Y=-7792 $D=0
M360 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=133735 $Y=-166 $D=0
M361 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=134095 $Y=-7792 $D=0
M362 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=134425 $Y=-166 $D=0
M363 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=134785 $Y=-7792 $D=0
M364 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=135115 $Y=-166 $D=0
M365 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=135475 $Y=-7792 $D=0
M366 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=135805 $Y=-166 $D=0
M367 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=136165 $Y=-7792 $D=0
M368 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=136495 $Y=-166 $D=0
M369 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=136855 $Y=-7792 $D=0
M370 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=137185 $Y=-166 $D=0
M371 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=137545 $Y=-7792 $D=0
M372 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=137875 $Y=-166 $D=0
M373 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=138235 $Y=-7792 $D=0
M374 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=138565 $Y=-166 $D=0
M375 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=138925 $Y=-7792 $D=0
M376 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=139255 $Y=-166 $D=0
M377 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=139615 $Y=-7792 $D=0
M378 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.425e-13 AS=1.275e-13 PD=5.7e-07 PS=5.1e-07 $X=139945 $Y=-166 $D=0
M379 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=140305 $Y=-7792 $D=0
M380 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.425e-13 PD=5.1e-07 PS=5.7e-07 $X=140695 $Y=-166 $D=0
M381 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=140995 $Y=-7792 $D=0
M382 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=141385 $Y=-166 $D=0
M383 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=141685 $Y=-7792 $D=0
M384 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=142075 $Y=-166 $D=0
M385 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=142375 $Y=-7792 $D=0
M386 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=142765 $Y=-166 $D=0
M387 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=143065 $Y=-7792 $D=0
M388 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=143455 $Y=-166 $D=0
M389 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=143755 $Y=-7792 $D=0
M390 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=144145 $Y=-166 $D=0
M391 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=144445 $Y=-7792 $D=0
M392 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=144835 $Y=-166 $D=0
M393 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=145135 $Y=-7792 $D=0
M394 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=145525 $Y=-166 $D=0
M395 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=145825 $Y=-7792 $D=0
M396 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=146215 $Y=-166 $D=0
M397 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=146515 $Y=-7792 $D=0
M398 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=146905 $Y=-166 $D=0
M399 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=147205 $Y=-7792 $D=0
M400 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=147595 $Y=-166 $D=0
M401 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=147895 $Y=-7792 $D=0
M402 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=148285 $Y=-166 $D=0
M403 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=148585 $Y=-7792 $D=0
M404 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=148975 $Y=-166 $D=0
M405 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=149275 $Y=-7792 $D=0
M406 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=149665 $Y=-166 $D=0
M407 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=149965 $Y=-7792 $D=0
M408 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=150355 $Y=-166 $D=0
M409 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=150655 $Y=-7792 $D=0
M410 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=151045 $Y=-166 $D=0
M411 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=151345 $Y=-7792 $D=0
M412 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=151735 $Y=-166 $D=0
M413 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=152035 $Y=-7792 $D=0
M414 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=152425 $Y=-166 $D=0
M415 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=152725 $Y=-7792 $D=0
M416 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=153115 $Y=-166 $D=0
M417 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=153415 $Y=-7792 $D=0
M418 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=153805 $Y=-166 $D=0
M419 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=154105 $Y=-7792 $D=0
M420 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=154495 $Y=-166 $D=0
M421 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=154795 $Y=-7792 $D=0
M422 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=155185 $Y=-166 $D=0
M423 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=155485 $Y=-7792 $D=0
M424 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=155875 $Y=-166 $D=0
M425 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=156175 $Y=-7792 $D=0
M426 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=156565 $Y=-166 $D=0
M427 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=156865 $Y=-7792 $D=0
M428 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=157255 $Y=-166 $D=0
M429 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=157555 $Y=-7792 $D=0
M430 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=157945 $Y=-166 $D=0
M431 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=158245 $Y=-7792 $D=0
M432 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=158635 $Y=-166 $D=0
M433 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=158935 $Y=-7792 $D=0
M434 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=159325 $Y=-166 $D=0
M435 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=159625 $Y=-7792 $D=0
M436 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=160015 $Y=-166 $D=0
M437 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=160315 $Y=-7792 $D=0
M438 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=160705 $Y=-166 $D=0
M439 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=161005 $Y=-7792 $D=0
M440 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=161395 $Y=-166 $D=0
M441 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=161695 $Y=-7792 $D=0
M442 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=162085 $Y=-166 $D=0
M443 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=162385 $Y=-7792 $D=0
M444 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=162775 $Y=-166 $D=0
M445 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=163075 $Y=-7792 $D=0
M446 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=163465 $Y=-166 $D=0
M447 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=163765 $Y=-7792 $D=0
M448 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=164155 $Y=-166 $D=0
M449 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=164455 $Y=-7792 $D=0
M450 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=164845 $Y=-166 $D=0
M451 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=165145 $Y=-7792 $D=0
M452 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=165535 $Y=-166 $D=0
M453 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=165835 $Y=-7792 $D=0
M454 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=166225 $Y=-166 $D=0
M455 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=166525 $Y=-7792 $D=0
M456 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=166915 $Y=-166 $D=0
M457 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=167215 $Y=-7792 $D=0
M458 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=167605 $Y=-166 $D=0
M459 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=167905 $Y=-7792 $D=0
M460 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=168295 $Y=-166 $D=0
M461 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=168595 $Y=-7792 $D=0
M462 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=168985 $Y=-166 $D=0
M463 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=169285 $Y=-7792 $D=0
M464 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=169675 $Y=-166 $D=0
M465 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=169975 $Y=-7792 $D=0
M466 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=170365 $Y=-166 $D=0
M467 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=170665 $Y=-7792 $D=0
M468 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=171055 $Y=-166 $D=0
M469 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=171355 $Y=-7792 $D=0
M470 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=171745 $Y=-166 $D=0
M471 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=172045 $Y=-7792 $D=0
M472 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=172435 $Y=-166 $D=0
M473 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=172735 $Y=-7792 $D=0
M474 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=173125 $Y=-166 $D=0
M475 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=173425 $Y=-7792 $D=0
M476 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=173815 $Y=-166 $D=0
M477 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=174115 $Y=-7792 $D=0
M478 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=174505 $Y=-166 $D=0
M479 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=174805 $Y=-7792 $D=0
M480 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=175195 $Y=-166 $D=0
M481 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=175495 $Y=-7792 $D=0
M482 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=175885 $Y=-166 $D=0
M483 17 16 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=176185 $Y=-7792 $D=0
M484 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=176575 $Y=-166 $D=0
M485 GND 16 17 GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=176875 $Y=-7792 $D=0
M486 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=177265 $Y=-166 $D=0
M487 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=177955 $Y=-166 $D=0
M488 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=178435 $Y=-7792 $D=0
M489 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=178645 $Y=-166 $D=0
M490 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=179125 $Y=-7792 $D=0
M491 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=179335 $Y=-166 $D=0
M492 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=179815 $Y=-7792 $D=0
M493 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=180025 $Y=-166 $D=0
M494 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=180505 $Y=-7792 $D=0
M495 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=180715 $Y=-166 $D=0
M496 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=181195 $Y=-7792 $D=0
M497 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=181405 $Y=-166 $D=0
M498 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=181885 $Y=-7792 $D=0
M499 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=182095 $Y=-166 $D=0
M500 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=182575 $Y=-7792 $D=0
M501 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=182785 $Y=-166 $D=0
M502 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=183265 $Y=-7792 $D=0
M503 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=183475 $Y=-166 $D=0
M504 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=183955 $Y=-7792 $D=0
M505 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=184165 $Y=-166 $D=0
M506 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=184645 $Y=-7792 $D=0
M507 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=184855 $Y=-166 $D=0
M508 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=185335 $Y=-7792 $D=0
M509 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=185545 $Y=-166 $D=0
M510 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=186025 $Y=-7792 $D=0
M511 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=186235 $Y=-166 $D=0
M512 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=186715 $Y=-7792 $D=0
M513 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=186925 $Y=-166 $D=0
M514 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=187405 $Y=-7792 $D=0
M515 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=187615 $Y=-166 $D=0
M516 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=188095 $Y=-7792 $D=0
M517 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=188305 $Y=-166 $D=0
M518 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=188785 $Y=-7792 $D=0
M519 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=188995 $Y=-166 $D=0
M520 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=189475 $Y=-7792 $D=0
M521 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=189685 $Y=-166 $D=0
M522 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=190165 $Y=-7792 $D=0
M523 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=190375 $Y=-166 $D=0
M524 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=190855 $Y=-7792 $D=0
M525 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=191065 $Y=-166 $D=0
M526 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=191545 $Y=-7792 $D=0
M527 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=191755 $Y=-166 $D=0
M528 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=192235 $Y=-7792 $D=0
M529 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=192445 $Y=-166 $D=0
M530 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=192925 $Y=-7792 $D=0
M531 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=193135 $Y=-166 $D=0
M532 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=193615 $Y=-7792 $D=0
M533 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=193825 $Y=-166 $D=0
M534 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=194305 $Y=-7792 $D=0
M535 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=194515 $Y=-166 $D=0
M536 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=194995 $Y=-7792 $D=0
M537 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=195205 $Y=-166 $D=0
M538 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=195685 $Y=-7792 $D=0
M539 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=195895 $Y=-166 $D=0
M540 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=196375 $Y=-7792 $D=0
M541 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=196585 $Y=-166 $D=0
M542 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=197065 $Y=-7792 $D=0
M543 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=197275 $Y=-166 $D=0
M544 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=197755 $Y=-7792 $D=0
M545 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=197965 $Y=-166 $D=0
M546 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=198445 $Y=-7792 $D=0
M547 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=198655 $Y=-166 $D=0
M548 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=199135 $Y=-7792 $D=0
M549 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=199345 $Y=-166 $D=0
M550 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=199825 $Y=-7792 $D=0
M551 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=200035 $Y=-166 $D=0
M552 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=200515 $Y=-7792 $D=0
M553 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=200725 $Y=-166 $D=0
M554 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=201205 $Y=-7792 $D=0
M555 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=201415 $Y=-166 $D=0
M556 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=201895 $Y=-7792 $D=0
M557 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=202105 $Y=-166 $D=0
M558 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=202585 $Y=-7792 $D=0
M559 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=202795 $Y=-166 $D=0
M560 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=203275 $Y=-7792 $D=0
M561 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=203485 $Y=-166 $D=0
M562 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=203965 $Y=-7792 $D=0
M563 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=204175 $Y=-166 $D=0
M564 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=204655 $Y=-7792 $D=0
M565 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=204865 $Y=-166 $D=0
M566 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=205345 $Y=-7792 $D=0
M567 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=205555 $Y=-166 $D=0
M568 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=206035 $Y=-7792 $D=0
M569 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=206245 $Y=-166 $D=0
M570 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=206725 $Y=-7792 $D=0
M571 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=206935 $Y=-166 $D=0
M572 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=207415 $Y=-7792 $D=0
M573 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=207625 $Y=-166 $D=0
M574 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=208105 $Y=-7792 $D=0
M575 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=208315 $Y=-166 $D=0
M576 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=208795 $Y=-7792 $D=0
M577 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=209005 $Y=-166 $D=0
M578 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=209485 $Y=-7792 $D=0
M579 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=209695 $Y=-166 $D=0
M580 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=210175 $Y=-7792 $D=0
M581 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=210385 $Y=-166 $D=0
M582 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=210865 $Y=-7792 $D=0
M583 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=211075 $Y=-166 $D=0
M584 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=211555 $Y=-7792 $D=0
M585 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=211765 $Y=-166 $D=0
M586 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=212245 $Y=-7792 $D=0
M587 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=212455 $Y=-166 $D=0
M588 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=212935 $Y=-7792 $D=0
M589 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=213145 $Y=-166 $D=0
M590 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=213625 $Y=-7792 $D=0
M591 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=213835 $Y=-166 $D=0
M592 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=214315 $Y=-7792 $D=0
M593 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=214525 $Y=-166 $D=0
M594 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=215005 $Y=-7792 $D=0
M595 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=215215 $Y=-166 $D=0
M596 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=215695 $Y=-7792 $D=0
M597 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=215905 $Y=-166 $D=0
M598 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=216385 $Y=-7792 $D=0
M599 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=216595 $Y=-166 $D=0
M600 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=217075 $Y=-7792 $D=0
M601 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=217285 $Y=-166 $D=0
M602 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=217765 $Y=-7792 $D=0
M603 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=217975 $Y=-166 $D=0
M604 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=218455 $Y=-7792 $D=0
M605 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=218665 $Y=-166 $D=0
M606 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=219145 $Y=-7792 $D=0
M607 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=219355 $Y=-166 $D=0
M608 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=219835 $Y=-7792 $D=0
M609 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=220045 $Y=-166 $D=0
M610 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=220525 $Y=-7792 $D=0
M611 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=220735 $Y=-166 $D=0
M612 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=221215 $Y=-7792 $D=0
M613 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=221425 $Y=-166 $D=0
M614 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=221905 $Y=-7792 $D=0
M615 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=222115 $Y=-166 $D=0
M616 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=222595 $Y=-7792 $D=0
M617 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=222805 $Y=-166 $D=0
M618 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=223285 $Y=-7792 $D=0
M619 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=223495 $Y=-166 $D=0
M620 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=223975 $Y=-7792 $D=0
M621 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=224185 $Y=-166 $D=0
M622 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=224665 $Y=-7792 $D=0
M623 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=224875 $Y=-166 $D=0
M624 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=225355 $Y=-7792 $D=0
M625 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=225565 $Y=-166 $D=0
M626 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=226045 $Y=-7792 $D=0
M627 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=226255 $Y=-166 $D=0
M628 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=226735 $Y=-7792 $D=0
M629 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=226945 $Y=-166 $D=0
M630 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=227425 $Y=-7792 $D=0
M631 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=227635 $Y=-166 $D=0
M632 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=228115 $Y=-7792 $D=0
M633 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=228325 $Y=-166 $D=0
M634 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=228805 $Y=-7792 $D=0
M635 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=229015 $Y=-166 $D=0
M636 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=229495 $Y=-7792 $D=0
M637 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=229705 $Y=-166 $D=0
M638 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=230185 $Y=-7792 $D=0
M639 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=230395 $Y=-166 $D=0
M640 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=230875 $Y=-7792 $D=0
M641 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=231085 $Y=-166 $D=0
M642 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=231565 $Y=-7792 $D=0
M643 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=231775 $Y=-166 $D=0
M644 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=232255 $Y=-7792 $D=0
M645 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=232465 $Y=-166 $D=0
M646 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=232945 $Y=-7792 $D=0
M647 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=233155 $Y=-166 $D=0
M648 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=233635 $Y=-7792 $D=0
M649 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=233845 $Y=-166 $D=0
M650 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=234325 $Y=-7792 $D=0
M651 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=234535 $Y=-166 $D=0
M652 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=235015 $Y=-7792 $D=0
M653 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=235225 $Y=-166 $D=0
M654 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=235705 $Y=-7792 $D=0
M655 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=235915 $Y=-166 $D=0
M656 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=236395 $Y=-7792 $D=0
M657 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=236605 $Y=-166 $D=0
M658 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=237085 $Y=-7792 $D=0
M659 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=237295 $Y=-166 $D=0
M660 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=237775 $Y=-7792 $D=0
M661 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=237985 $Y=-166 $D=0
M662 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=238465 $Y=-7792 $D=0
M663 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=238675 $Y=-166 $D=0
M664 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=239155 $Y=-7792 $D=0
M665 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=239365 $Y=-166 $D=0
M666 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.425e-13 AS=1.275e-13 PD=5.7e-07 PS=5.1e-07 $X=239845 $Y=-7792 $D=0
M667 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=240055 $Y=-166 $D=0
M668 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.425e-13 PD=5.1e-07 PS=5.7e-07 $X=240595 $Y=-7792 $D=0
M669 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=240745 $Y=-166 $D=0
M670 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=241285 $Y=-7792 $D=0
M671 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=241435 $Y=-166 $D=0
M672 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=241975 $Y=-7792 $D=0
M673 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=242125 $Y=-166 $D=0
M674 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=242665 $Y=-7792 $D=0
M675 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=242815 $Y=-166 $D=0
M676 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=243355 $Y=-7792 $D=0
M677 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=243505 $Y=-166 $D=0
M678 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=244045 $Y=-7792 $D=0
M679 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=244195 $Y=-166 $D=0
M680 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=244735 $Y=-7792 $D=0
M681 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=244885 $Y=-166 $D=0
M682 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=245425 $Y=-7792 $D=0
M683 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=245575 $Y=-166 $D=0
M684 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=246115 $Y=-7792 $D=0
M685 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=246265 $Y=-166 $D=0
M686 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=246805 $Y=-7792 $D=0
M687 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=246955 $Y=-166 $D=0
M688 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=247495 $Y=-7792 $D=0
M689 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=247645 $Y=-166 $D=0
M690 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=248185 $Y=-7792 $D=0
M691 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=248335 $Y=-166 $D=0
M692 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=248875 $Y=-7792 $D=0
M693 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=249025 $Y=-166 $D=0
M694 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=249565 $Y=-7792 $D=0
M695 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=249715 $Y=-166 $D=0
M696 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=250255 $Y=-7792 $D=0
M697 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=250405 $Y=-166 $D=0
M698 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=250945 $Y=-7792 $D=0
M699 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=251095 $Y=-166 $D=0
M700 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=251635 $Y=-7792 $D=0
M701 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=251785 $Y=-166 $D=0
M702 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=252325 $Y=-7792 $D=0
M703 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=252475 $Y=-166 $D=0
M704 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=253015 $Y=-7792 $D=0
M705 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=253165 $Y=-166 $D=0
M706 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=253705 $Y=-7792 $D=0
M707 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=253855 $Y=-166 $D=0
M708 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=254395 $Y=-7792 $D=0
M709 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=254545 $Y=-166 $D=0
M710 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=255085 $Y=-7792 $D=0
M711 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=255235 $Y=-166 $D=0
M712 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=255775 $Y=-7792 $D=0
M713 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=255925 $Y=-166 $D=0
M714 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=256465 $Y=-7792 $D=0
M715 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=256615 $Y=-166 $D=0
M716 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=257155 $Y=-7792 $D=0
M717 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=257305 $Y=-166 $D=0
M718 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=257845 $Y=-7792 $D=0
M719 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=257995 $Y=-166 $D=0
M720 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=258535 $Y=-7792 $D=0
M721 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=258685 $Y=-166 $D=0
M722 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=259225 $Y=-7792 $D=0
M723 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=259375 $Y=-166 $D=0
M724 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=259915 $Y=-7792 $D=0
M725 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=260065 $Y=-166 $D=0
M726 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=260605 $Y=-7792 $D=0
M727 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=260755 $Y=-166 $D=0
M728 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=261295 $Y=-7792 $D=0
M729 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=261445 $Y=-166 $D=0
M730 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=261985 $Y=-7792 $D=0
M731 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=262135 $Y=-166 $D=0
M732 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=262675 $Y=-7792 $D=0
M733 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=262825 $Y=-166 $D=0
M734 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=263365 $Y=-7792 $D=0
M735 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=263515 $Y=-166 $D=0
M736 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=264055 $Y=-7792 $D=0
M737 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=264205 $Y=-166 $D=0
M738 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=264745 $Y=-7792 $D=0
M739 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=264895 $Y=-166 $D=0
M740 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=265435 $Y=-7792 $D=0
M741 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=265585 $Y=-166 $D=0
M742 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=266125 $Y=-7792 $D=0
M743 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=266275 $Y=-166 $D=0
M744 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=266815 $Y=-7792 $D=0
M745 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=266965 $Y=-166 $D=0
M746 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=267505 $Y=-7792 $D=0
M747 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=267655 $Y=-166 $D=0
M748 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=268195 $Y=-7792 $D=0
M749 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=268345 $Y=-166 $D=0
M750 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=268885 $Y=-7792 $D=0
M751 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=269035 $Y=-166 $D=0
M752 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=269575 $Y=-7792 $D=0
M753 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=269725 $Y=-166 $D=0
M754 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=270265 $Y=-7792 $D=0
M755 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=270415 $Y=-166 $D=0
M756 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=270955 $Y=-7792 $D=0
M757 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=271105 $Y=-166 $D=0
M758 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=271645 $Y=-7792 $D=0
M759 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=271795 $Y=-166 $D=0
M760 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=272335 $Y=-7792 $D=0
M761 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=272485 $Y=-166 $D=0
M762 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=273025 $Y=-7792 $D=0
M763 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=273175 $Y=-166 $D=0
M764 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=273715 $Y=-7792 $D=0
M765 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=273865 $Y=-166 $D=0
M766 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=274405 $Y=-7792 $D=0
M767 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=274555 $Y=-166 $D=0
M768 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=275095 $Y=-7792 $D=0
M769 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=275245 $Y=-166 $D=0
M770 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=275785 $Y=-7792 $D=0
M771 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=275935 $Y=-166 $D=0
M772 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=276475 $Y=-7792 $D=0
M773 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=276625 $Y=-166 $D=0
M774 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=277165 $Y=-7792 $D=0
M775 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=277315 $Y=-166 $D=0
M776 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=277855 $Y=-7792 $D=0
M777 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=278005 $Y=-166 $D=0
M778 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=278545 $Y=-7792 $D=0
M779 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=278695 $Y=-166 $D=0
M780 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=279235 $Y=-7792 $D=0
M781 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=279385 $Y=-166 $D=0
M782 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=279925 $Y=-7792 $D=0
M783 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=280075 $Y=-166 $D=0
M784 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=280615 $Y=-7792 $D=0
M785 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=280765 $Y=-166 $D=0
M786 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=281305 $Y=-7792 $D=0
M787 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=281455 $Y=-166 $D=0
M788 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=281995 $Y=-7792 $D=0
M789 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=282145 $Y=-166 $D=0
M790 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=282685 $Y=-7792 $D=0
M791 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=282835 $Y=-166 $D=0
M792 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=283375 $Y=-7792 $D=0
M793 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=283525 $Y=-166 $D=0
M794 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=284065 $Y=-7792 $D=0
M795 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=284215 $Y=-166 $D=0
M796 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=284755 $Y=-7792 $D=0
M797 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=284905 $Y=-166 $D=0
M798 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=285445 $Y=-7792 $D=0
M799 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=285595 $Y=-166 $D=0
M800 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=286135 $Y=-7792 $D=0
M801 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=286285 $Y=-166 $D=0
M802 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=286825 $Y=-7792 $D=0
M803 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=286975 $Y=-166 $D=0
M804 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=287515 $Y=-7792 $D=0
M805 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=287665 $Y=-166 $D=0
M806 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=288205 $Y=-7792 $D=0
M807 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=288355 $Y=-166 $D=0
M808 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=288895 $Y=-7792 $D=0
M809 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=289045 $Y=-166 $D=0
M810 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=289585 $Y=-7792 $D=0
M811 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=289735 $Y=-166 $D=0
M812 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=290275 $Y=-7792 $D=0
M813 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=290425 $Y=-166 $D=0
M814 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=290965 $Y=-7792 $D=0
M815 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=291115 $Y=-166 $D=0
M816 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=291655 $Y=-7792 $D=0
M817 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=291805 $Y=-166 $D=0
M818 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=292345 $Y=-7792 $D=0
M819 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=292495 $Y=-166 $D=0
M820 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=293035 $Y=-7792 $D=0
M821 GND 15 Vbout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=293185 $Y=-166 $D=0
M822 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=293725 $Y=-7792 $D=0
M823 Vbout 15 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=293875 $Y=-166 $D=0
M824 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=294415 $Y=-7792 $D=0
M825 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=295105 $Y=-7792 $D=0
M826 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=295795 $Y=-7792 $D=0
M827 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=296485 $Y=-7792 $D=0
M828 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=297175 $Y=-7792 $D=0
M829 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=297865 $Y=-7792 $D=0
M830 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=298555 $Y=-7792 $D=0
M831 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=299245 $Y=-7792 $D=0
M832 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=299935 $Y=-7792 $D=0
M833 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=300625 $Y=-7792 $D=0
M834 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=301315 $Y=-7792 $D=0
M835 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=302005 $Y=-7792 $D=0
M836 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=302695 $Y=-7792 $D=0
M837 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=303385 $Y=-7792 $D=0
M838 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=304075 $Y=-7792 $D=0
M839 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=304765 $Y=-7792 $D=0
M840 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=305455 $Y=-7792 $D=0
M841 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=306145 $Y=-7792 $D=0
M842 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=306835 $Y=-7792 $D=0
M843 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=307525 $Y=-7792 $D=0
M844 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=308215 $Y=-7792 $D=0
M845 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=308905 $Y=-7792 $D=0
M846 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=309595 $Y=-7792 $D=0
M847 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=310285 $Y=-7792 $D=0
M848 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=310975 $Y=-7792 $D=0
M849 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=311665 $Y=-7792 $D=0
M850 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=312355 $Y=-7792 $D=0
M851 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=313045 $Y=-7792 $D=0
M852 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=313735 $Y=-7792 $D=0
M853 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=314425 $Y=-7792 $D=0
M854 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=315115 $Y=-7792 $D=0
M855 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=315805 $Y=-7792 $D=0
M856 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=316495 $Y=-7792 $D=0
M857 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=317185 $Y=-7792 $D=0
M858 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=317875 $Y=-7792 $D=0
M859 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=318565 $Y=-7792 $D=0
M860 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=319255 $Y=-7792 $D=0
M861 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=319945 $Y=-7792 $D=0
M862 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=320635 $Y=-7792 $D=0
M863 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=321325 $Y=-7792 $D=0
M864 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=322015 $Y=-7792 $D=0
M865 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=322705 $Y=-7792 $D=0
M866 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=323395 $Y=-7792 $D=0
M867 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=324085 $Y=-7792 $D=0
M868 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=324775 $Y=-7792 $D=0
M869 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=325465 $Y=-7792 $D=0
M870 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=326155 $Y=-7792 $D=0
M871 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=326845 $Y=-7792 $D=0
M872 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=327535 $Y=-7792 $D=0
M873 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=328225 $Y=-7792 $D=0
M874 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=328915 $Y=-7792 $D=0
M875 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=329605 $Y=-7792 $D=0
M876 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=330295 $Y=-7792 $D=0
M877 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=330985 $Y=-7792 $D=0
M878 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=331675 $Y=-7792 $D=0
M879 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=332365 $Y=-7792 $D=0
M880 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=333055 $Y=-7792 $D=0
M881 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=333745 $Y=-7792 $D=0
M882 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=334435 $Y=-7792 $D=0
M883 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=335125 $Y=-7792 $D=0
M884 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=335815 $Y=-7792 $D=0
M885 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=336505 $Y=-7792 $D=0
M886 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=337195 $Y=-7792 $D=0
M887 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=337885 $Y=-7792 $D=0
M888 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=338575 $Y=-7792 $D=0
M889 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=339265 $Y=-7792 $D=0
M890 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=339955 $Y=-7792 $D=0
M891 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=340645 $Y=-7792 $D=0
M892 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=341335 $Y=-7792 $D=0
M893 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=342025 $Y=-7792 $D=0
M894 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=342715 $Y=-7792 $D=0
M895 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=343405 $Y=-7792 $D=0
M896 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=344095 $Y=-7792 $D=0
M897 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=344785 $Y=-7792 $D=0
M898 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=345475 $Y=-7792 $D=0
M899 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=346165 $Y=-7792 $D=0
M900 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=346855 $Y=-7792 $D=0
M901 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=347545 $Y=-7792 $D=0
M902 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=348235 $Y=-7792 $D=0
M903 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=348925 $Y=-7792 $D=0
M904 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=349615 $Y=-7792 $D=0
M905 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=350305 $Y=-7792 $D=0
M906 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=350995 $Y=-7792 $D=0
M907 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=351685 $Y=-7792 $D=0
M908 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=352375 $Y=-7792 $D=0
M909 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=353065 $Y=-7792 $D=0
M910 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=353755 $Y=-7792 $D=0
M911 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=354445 $Y=-7792 $D=0
M912 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=355135 $Y=-7792 $D=0
M913 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=355825 $Y=-7792 $D=0
M914 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=356515 $Y=-7792 $D=0
M915 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=357205 $Y=-7792 $D=0
M916 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=357895 $Y=-7792 $D=0
M917 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=358585 $Y=-7792 $D=0
M918 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=359275 $Y=-7792 $D=0
M919 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=359965 $Y=-7792 $D=0
M920 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=360655 $Y=-7792 $D=0
M921 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=361345 $Y=-7792 $D=0
M922 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=362035 $Y=-7792 $D=0
M923 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=362725 $Y=-7792 $D=0
M924 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=363415 $Y=-7792 $D=0
M925 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=364105 $Y=-7792 $D=0
M926 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=364795 $Y=-7792 $D=0
M927 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=365485 $Y=-7792 $D=0
M928 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=366175 $Y=-7792 $D=0
M929 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=366865 $Y=-7792 $D=0
M930 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=367555 $Y=-7792 $D=0
M931 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=368245 $Y=-7792 $D=0
M932 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=368935 $Y=-7792 $D=0
M933 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=369625 $Y=-7792 $D=0
M934 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=370315 $Y=-7792 $D=0
M935 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=371005 $Y=-7792 $D=0
M936 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=371695 $Y=-7792 $D=0
M937 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=372385 $Y=-7792 $D=0
M938 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=373075 $Y=-7792 $D=0
M939 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=373765 $Y=-7792 $D=0
M940 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=374455 $Y=-7792 $D=0
M941 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=375145 $Y=-7792 $D=0
M942 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=375835 $Y=-7792 $D=0
M943 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=376525 $Y=-7792 $D=0
M944 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=377215 $Y=-7792 $D=0
M945 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=377905 $Y=-7792 $D=0
M946 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=378595 $Y=-7792 $D=0
M947 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=379285 $Y=-7792 $D=0
M948 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=379975 $Y=-7792 $D=0
M949 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=380665 $Y=-7792 $D=0
M950 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=381355 $Y=-7792 $D=0
M951 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=382045 $Y=-7792 $D=0
M952 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=382735 $Y=-7792 $D=0
M953 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=383425 $Y=-7792 $D=0
M954 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=384115 $Y=-7792 $D=0
M955 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=384805 $Y=-7792 $D=0
M956 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=385495 $Y=-7792 $D=0
M957 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=386185 $Y=-7792 $D=0
M958 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=386875 $Y=-7792 $D=0
M959 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=387565 $Y=-7792 $D=0
M960 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=388255 $Y=-7792 $D=0
M961 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=388945 $Y=-7792 $D=0
M962 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=389635 $Y=-7792 $D=0
M963 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=390325 $Y=-7792 $D=0
M964 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=391015 $Y=-7792 $D=0
M965 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=391705 $Y=-7792 $D=0
M966 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=392395 $Y=-7792 $D=0
M967 GND 17 19 GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=393085 $Y=-7792 $D=0
M968 19 17 GND GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=393775 $Y=-7792 $D=0
M969 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=2.45e-13 PD=5.1e-07 PS=1.48e-06 $X=395335 $Y=-7792 $D=0
M970 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=396025 $Y=-7792 $D=0
M971 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=396715 $Y=-7792 $D=0
M972 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=397405 $Y=-7792 $D=0
M973 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=398095 $Y=-7792 $D=0
M974 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=398785 $Y=-7792 $D=0
M975 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=399475 $Y=-7792 $D=0
M976 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=400165 $Y=-7792 $D=0
M977 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=400855 $Y=-7792 $D=0
M978 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=401545 $Y=-7792 $D=0
M979 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=402235 $Y=-7792 $D=0
M980 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=402925 $Y=-7792 $D=0
M981 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=403615 $Y=-7792 $D=0
M982 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=404305 $Y=-7792 $D=0
M983 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=404995 $Y=-7792 $D=0
M984 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=405685 $Y=-7792 $D=0
M985 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=406375 $Y=-7792 $D=0
M986 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=407065 $Y=-7792 $D=0
M987 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=407755 $Y=-7792 $D=0
M988 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=408445 $Y=-7792 $D=0
M989 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=409135 $Y=-7792 $D=0
M990 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=409825 $Y=-7792 $D=0
M991 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=410515 $Y=-7792 $D=0
M992 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=411205 $Y=-7792 $D=0
M993 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=411895 $Y=-7792 $D=0
M994 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=412585 $Y=-7792 $D=0
M995 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=413275 $Y=-7792 $D=0
M996 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=413965 $Y=-7792 $D=0
M997 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=414655 $Y=-7792 $D=0
M998 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=415345 $Y=-7792 $D=0
M999 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=416035 $Y=-7792 $D=0
M1000 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=416725 $Y=-7792 $D=0
M1001 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=417415 $Y=-7792 $D=0
M1002 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=418105 $Y=-7792 $D=0
M1003 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=418795 $Y=-7792 $D=0
M1004 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=419485 $Y=-7792 $D=0
M1005 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=420175 $Y=-7792 $D=0
M1006 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=420865 $Y=-7792 $D=0
M1007 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=421555 $Y=-7792 $D=0
M1008 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=422245 $Y=-7792 $D=0
M1009 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=422935 $Y=-7792 $D=0
M1010 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=423625 $Y=-7792 $D=0
M1011 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=424315 $Y=-7792 $D=0
M1012 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=425005 $Y=-7792 $D=0
M1013 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=425695 $Y=-7792 $D=0
M1014 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=426385 $Y=-7792 $D=0
M1015 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=427075 $Y=-7792 $D=0
M1016 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=427765 $Y=-7792 $D=0
M1017 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=428455 $Y=-7792 $D=0
M1018 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=429145 $Y=-7792 $D=0
M1019 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=429835 $Y=-7792 $D=0
M1020 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=430525 $Y=-7792 $D=0
M1021 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=431215 $Y=-7792 $D=0
M1022 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=431905 $Y=-7792 $D=0
M1023 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=432595 $Y=-7792 $D=0
M1024 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=433285 $Y=-7792 $D=0
M1025 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=433975 $Y=-7792 $D=0
M1026 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=434665 $Y=-7792 $D=0
M1027 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=435355 $Y=-7792 $D=0
M1028 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=436045 $Y=-7792 $D=0
M1029 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=436735 $Y=-7792 $D=0
M1030 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=437425 $Y=-7792 $D=0
M1031 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=438115 $Y=-7792 $D=0
M1032 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=438805 $Y=-7792 $D=0
M1033 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=439495 $Y=-7792 $D=0
M1034 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=440185 $Y=-7792 $D=0
M1035 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=440875 $Y=-7792 $D=0
M1036 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=441565 $Y=-7792 $D=0
M1037 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=442255 $Y=-7792 $D=0
M1038 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=442945 $Y=-7792 $D=0
M1039 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=443635 $Y=-7792 $D=0
M1040 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=444325 $Y=-7792 $D=0
M1041 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=445015 $Y=-7792 $D=0
M1042 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=445705 $Y=-7792 $D=0
M1043 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=446395 $Y=-7792 $D=0
M1044 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=447085 $Y=-7792 $D=0
M1045 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=447775 $Y=-7792 $D=0
M1046 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=448465 $Y=-7792 $D=0
M1047 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=449155 $Y=-7792 $D=0
M1048 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=449845 $Y=-7792 $D=0
M1049 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=450535 $Y=-7792 $D=0
M1050 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=451225 $Y=-7792 $D=0
M1051 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=451915 $Y=-7792 $D=0
M1052 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=452605 $Y=-7792 $D=0
M1053 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=453295 $Y=-7792 $D=0
M1054 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=453985 $Y=-7792 $D=0
M1055 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=454675 $Y=-7792 $D=0
M1056 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=455365 $Y=-7792 $D=0
M1057 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=456055 $Y=-7792 $D=0
M1058 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.425e-13 AS=1.275e-13 PD=5.7e-07 PS=5.1e-07 $X=456745 $Y=-7792 $D=0
M1059 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.425e-13 PD=5.1e-07 PS=5.7e-07 $X=457495 $Y=-7792 $D=0
M1060 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=458185 $Y=-7792 $D=0
M1061 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=458875 $Y=-7792 $D=0
M1062 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=459565 $Y=-7792 $D=0
M1063 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=460255 $Y=-7792 $D=0
M1064 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=460945 $Y=-7792 $D=0
M1065 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=461635 $Y=-7792 $D=0
M1066 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=462325 $Y=-7792 $D=0
M1067 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=463015 $Y=-7792 $D=0
M1068 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=463705 $Y=-7792 $D=0
M1069 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=464395 $Y=-7792 $D=0
M1070 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=465085 $Y=-7792 $D=0
M1071 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=465775 $Y=-7792 $D=0
M1072 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=466465 $Y=-7792 $D=0
M1073 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=467155 $Y=-7792 $D=0
M1074 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=467845 $Y=-7792 $D=0
M1075 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=468535 $Y=-7792 $D=0
M1076 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=469225 $Y=-7792 $D=0
M1077 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=469915 $Y=-7792 $D=0
M1078 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=470605 $Y=-7792 $D=0
M1079 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=471295 $Y=-7792 $D=0
M1080 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=471985 $Y=-7792 $D=0
M1081 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=472675 $Y=-7792 $D=0
M1082 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=473365 $Y=-7792 $D=0
M1083 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=474055 $Y=-7792 $D=0
M1084 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=474745 $Y=-7792 $D=0
M1085 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=475435 $Y=-7792 $D=0
M1086 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=476125 $Y=-7792 $D=0
M1087 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=476815 $Y=-7792 $D=0
M1088 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=477505 $Y=-7792 $D=0
M1089 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=478195 $Y=-7792 $D=0
M1090 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=478885 $Y=-7792 $D=0
M1091 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=479575 $Y=-7792 $D=0
M1092 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=480265 $Y=-7792 $D=0
M1093 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=480955 $Y=-7792 $D=0
M1094 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=481645 $Y=-7792 $D=0
M1095 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=482335 $Y=-7792 $D=0
M1096 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=483025 $Y=-7792 $D=0
M1097 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=483715 $Y=-7792 $D=0
M1098 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=484405 $Y=-7792 $D=0
M1099 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=485095 $Y=-7792 $D=0
M1100 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=485785 $Y=-7792 $D=0
M1101 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=486475 $Y=-7792 $D=0
M1102 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=487165 $Y=-7792 $D=0
M1103 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=487855 $Y=-7792 $D=0
M1104 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=488545 $Y=-7792 $D=0
M1105 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=489235 $Y=-7792 $D=0
M1106 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=489925 $Y=-7792 $D=0
M1107 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=490615 $Y=-7792 $D=0
M1108 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=491305 $Y=-7792 $D=0
M1109 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=491995 $Y=-7792 $D=0
M1110 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=492685 $Y=-7792 $D=0
M1111 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=493375 $Y=-7792 $D=0
M1112 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=494065 $Y=-7792 $D=0
M1113 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=494755 $Y=-7792 $D=0
M1114 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=495445 $Y=-7792 $D=0
M1115 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=496135 $Y=-7792 $D=0
M1116 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=496825 $Y=-7792 $D=0
M1117 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=497515 $Y=-7792 $D=0
M1118 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=498205 $Y=-7792 $D=0
M1119 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=498895 $Y=-7792 $D=0
M1120 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=499585 $Y=-7792 $D=0
M1121 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=500275 $Y=-7792 $D=0
M1122 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=500965 $Y=-7792 $D=0
M1123 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=501655 $Y=-7792 $D=0
M1124 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=502345 $Y=-7792 $D=0
M1125 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=503035 $Y=-7792 $D=0
M1126 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=503725 $Y=-7792 $D=0
M1127 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=504415 $Y=-7792 $D=0
M1128 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=505105 $Y=-7792 $D=0
M1129 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=505795 $Y=-7792 $D=0
M1130 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=506485 $Y=-7792 $D=0
M1131 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=507175 $Y=-7792 $D=0
M1132 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=507865 $Y=-7792 $D=0
M1133 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=508555 $Y=-7792 $D=0
M1134 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=509245 $Y=-7792 $D=0
M1135 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=509935 $Y=-7792 $D=0
M1136 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=510625 $Y=-7792 $D=0
M1137 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=511315 $Y=-7792 $D=0
M1138 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=512005 $Y=-7792 $D=0
M1139 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=512695 $Y=-7792 $D=0
M1140 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=513385 $Y=-7792 $D=0
M1141 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=514075 $Y=-7792 $D=0
M1142 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=514765 $Y=-7792 $D=0
M1143 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=515455 $Y=-7792 $D=0
M1144 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=516145 $Y=-7792 $D=0
M1145 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=516835 $Y=-7792 $D=0
M1146 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=517525 $Y=-7792 $D=0
M1147 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=518215 $Y=-7792 $D=0
M1148 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=518905 $Y=-7792 $D=0
M1149 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=519595 $Y=-7792 $D=0
M1150 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=520285 $Y=-7792 $D=0
M1151 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=520975 $Y=-7792 $D=0
M1152 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=521665 $Y=-7792 $D=0
M1153 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=522355 $Y=-7792 $D=0
M1154 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=523045 $Y=-7792 $D=0
M1155 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=523735 $Y=-7792 $D=0
M1156 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=524425 $Y=-7792 $D=0
M1157 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=525115 $Y=-7792 $D=0
M1158 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=525805 $Y=-7792 $D=0
M1159 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=526495 $Y=-7792 $D=0
M1160 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=527185 $Y=-7792 $D=0
M1161 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=527875 $Y=-7792 $D=0
M1162 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=528565 $Y=-7792 $D=0
M1163 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=529255 $Y=-7792 $D=0
M1164 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=529945 $Y=-7792 $D=0
M1165 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=530635 $Y=-7792 $D=0
M1166 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=531325 $Y=-7792 $D=0
M1167 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=532015 $Y=-7792 $D=0
M1168 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=532705 $Y=-7792 $D=0
M1169 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=533395 $Y=-7792 $D=0
M1170 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=534085 $Y=-7792 $D=0
M1171 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=534775 $Y=-7792 $D=0
M1172 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=535465 $Y=-7792 $D=0
M1173 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=536155 $Y=-7792 $D=0
M1174 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=536845 $Y=-7792 $D=0
M1175 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=537535 $Y=-7792 $D=0
M1176 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=538225 $Y=-7792 $D=0
M1177 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=538915 $Y=-7792 $D=0
M1178 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=539605 $Y=-7792 $D=0
M1179 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=540295 $Y=-7792 $D=0
M1180 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=540985 $Y=-7792 $D=0
M1181 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=541675 $Y=-7792 $D=0
M1182 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=542365 $Y=-7792 $D=0
M1183 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=543055 $Y=-7792 $D=0
M1184 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=543745 $Y=-7792 $D=0
M1185 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=544435 $Y=-7792 $D=0
M1186 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=545125 $Y=-7792 $D=0
M1187 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=545815 $Y=-7792 $D=0
M1188 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=546505 $Y=-7792 $D=0
M1189 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=547195 $Y=-7792 $D=0
M1190 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=547885 $Y=-7792 $D=0
M1191 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=548575 $Y=-7792 $D=0
M1192 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=549265 $Y=-7792 $D=0
M1193 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=549955 $Y=-7792 $D=0
M1194 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=550645 $Y=-7792 $D=0
M1195 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=551335 $Y=-7792 $D=0
M1196 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=552025 $Y=-7792 $D=0
M1197 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=552715 $Y=-7792 $D=0
M1198 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=553405 $Y=-7792 $D=0
M1199 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=554095 $Y=-7792 $D=0
M1200 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=554785 $Y=-7792 $D=0
M1201 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=555475 $Y=-7792 $D=0
M1202 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=556165 $Y=-7792 $D=0
M1203 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=556855 $Y=-7792 $D=0
M1204 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=557545 $Y=-7792 $D=0
M1205 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=558235 $Y=-7792 $D=0
M1206 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=558925 $Y=-7792 $D=0
M1207 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=559615 $Y=-7792 $D=0
M1208 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=560305 $Y=-7792 $D=0
M1209 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=560995 $Y=-7792 $D=0
M1210 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=561685 $Y=-7792 $D=0
M1211 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=562375 $Y=-7792 $D=0
M1212 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=563065 $Y=-7792 $D=0
M1213 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=563755 $Y=-7792 $D=0
M1214 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=564445 $Y=-7792 $D=0
M1215 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=565135 $Y=-7792 $D=0
M1216 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=565825 $Y=-7792 $D=0
M1217 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=566515 $Y=-7792 $D=0
M1218 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=567205 $Y=-7792 $D=0
M1219 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=567895 $Y=-7792 $D=0
M1220 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=568585 $Y=-7792 $D=0
M1221 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=569275 $Y=-7792 $D=0
M1222 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=569965 $Y=-7792 $D=0
M1223 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=570655 $Y=-7792 $D=0
M1224 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=571345 $Y=-7792 $D=0
M1225 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=572035 $Y=-7792 $D=0
M1226 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=572725 $Y=-7792 $D=0
M1227 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=573415 $Y=-7792 $D=0
M1228 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=574105 $Y=-7792 $D=0
M1229 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=574795 $Y=-7792 $D=0
M1230 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=575485 $Y=-7792 $D=0
M1231 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=576175 $Y=-7792 $D=0
M1232 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=576865 $Y=-7792 $D=0
M1233 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=577555 $Y=-7792 $D=0
M1234 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=578245 $Y=-7792 $D=0
M1235 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=578935 $Y=-7792 $D=0
M1236 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=579625 $Y=-7792 $D=0
M1237 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=580315 $Y=-7792 $D=0
M1238 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=581005 $Y=-7792 $D=0
M1239 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=581695 $Y=-7792 $D=0
M1240 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=582385 $Y=-7792 $D=0
M1241 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=583075 $Y=-7792 $D=0
M1242 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=583765 $Y=-7792 $D=0
M1243 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=584455 $Y=-7792 $D=0
M1244 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=585145 $Y=-7792 $D=0
M1245 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=585835 $Y=-7792 $D=0
M1246 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=586525 $Y=-7792 $D=0
M1247 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=587215 $Y=-7792 $D=0
M1248 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=587905 $Y=-7792 $D=0
M1249 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=588595 $Y=-7792 $D=0
M1250 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=589285 $Y=-7792 $D=0
M1251 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=589975 $Y=-7792 $D=0
M1252 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=590665 $Y=-7792 $D=0
M1253 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=591355 $Y=-7792 $D=0
M1254 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=592045 $Y=-7792 $D=0
M1255 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=592735 $Y=-7792 $D=0
M1256 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=593425 $Y=-7792 $D=0
M1257 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=594115 $Y=-7792 $D=0
M1258 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=594805 $Y=-7792 $D=0
M1259 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=595495 $Y=-7792 $D=0
M1260 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=596185 $Y=-7792 $D=0
M1261 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=596875 $Y=-7792 $D=0
M1262 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=597565 $Y=-7792 $D=0
M1263 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=598255 $Y=-7792 $D=0
M1264 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=598945 $Y=-7792 $D=0
M1265 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=599635 $Y=-7792 $D=0
M1266 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=600325 $Y=-7792 $D=0
M1267 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=601015 $Y=-7792 $D=0
M1268 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=601705 $Y=-7792 $D=0
M1269 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=602395 $Y=-7792 $D=0
M1270 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=603085 $Y=-7792 $D=0
M1271 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=603775 $Y=-7792 $D=0
M1272 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=604465 $Y=-7792 $D=0
M1273 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=605155 $Y=-7792 $D=0
M1274 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=605845 $Y=-7792 $D=0
M1275 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=606535 $Y=-7792 $D=0
M1276 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=607225 $Y=-7792 $D=0
M1277 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=607915 $Y=-7792 $D=0
M1278 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=608605 $Y=-7792 $D=0
M1279 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=609295 $Y=-7792 $D=0
M1280 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=609985 $Y=-7792 $D=0
M1281 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=610675 $Y=-7792 $D=0
M1282 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=611365 $Y=-7792 $D=0
M1283 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=612055 $Y=-7792 $D=0
M1284 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=612745 $Y=-7792 $D=0
M1285 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=613435 $Y=-7792 $D=0
M1286 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=614125 $Y=-7792 $D=0
M1287 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=614815 $Y=-7792 $D=0
M1288 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=615505 $Y=-7792 $D=0
M1289 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=616195 $Y=-7792 $D=0
M1290 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=616885 $Y=-7792 $D=0
M1291 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=617575 $Y=-7792 $D=0
M1292 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=618265 $Y=-7792 $D=0
M1293 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=618955 $Y=-7792 $D=0
M1294 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=619645 $Y=-7792 $D=0
M1295 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=620335 $Y=-7792 $D=0
M1296 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=621025 $Y=-7792 $D=0
M1297 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=621715 $Y=-7792 $D=0
M1298 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=622405 $Y=-7792 $D=0
M1299 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=623095 $Y=-7792 $D=0
M1300 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=623785 $Y=-7792 $D=0
M1301 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=624475 $Y=-7792 $D=0
M1302 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=625165 $Y=-7792 $D=0
M1303 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=625855 $Y=-7792 $D=0
M1304 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=626545 $Y=-7792 $D=0
M1305 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=627235 $Y=-7792 $D=0
M1306 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=627925 $Y=-7792 $D=0
M1307 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=628615 $Y=-7792 $D=0
M1308 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=629305 $Y=-7792 $D=0
M1309 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=629995 $Y=-7792 $D=0
M1310 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=630685 $Y=-7792 $D=0
M1311 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=631375 $Y=-7792 $D=0
M1312 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=632065 $Y=-7792 $D=0
M1313 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=632755 $Y=-7792 $D=0
M1314 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=633445 $Y=-7792 $D=0
M1315 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=634135 $Y=-7792 $D=0
M1316 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=634825 $Y=-7792 $D=0
M1317 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=635515 $Y=-7792 $D=0
M1318 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=636205 $Y=-7792 $D=0
M1319 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=636895 $Y=-7792 $D=0
M1320 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=637585 $Y=-7792 $D=0
M1321 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=638275 $Y=-7792 $D=0
M1322 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=638965 $Y=-7792 $D=0
M1323 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=639655 $Y=-7792 $D=0
M1324 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=640345 $Y=-7792 $D=0
M1325 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=641035 $Y=-7792 $D=0
M1326 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=641725 $Y=-7792 $D=0
M1327 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=642415 $Y=-7792 $D=0
M1328 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=643105 $Y=-7792 $D=0
M1329 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=643795 $Y=-7792 $D=0
M1330 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=644485 $Y=-7792 $D=0
M1331 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=645175 $Y=-7792 $D=0
M1332 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=645865 $Y=-7792 $D=0
M1333 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=646555 $Y=-7792 $D=0
M1334 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=647245 $Y=-7792 $D=0
M1335 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=647935 $Y=-7792 $D=0
M1336 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=648625 $Y=-7792 $D=0
M1337 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=649315 $Y=-7792 $D=0
M1338 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=650005 $Y=-7792 $D=0
M1339 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=650695 $Y=-7792 $D=0
M1340 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=651385 $Y=-7792 $D=0
M1341 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=652075 $Y=-7792 $D=0
M1342 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=652765 $Y=-7792 $D=0
M1343 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=653455 $Y=-7792 $D=0
M1344 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=654145 $Y=-7792 $D=0
M1345 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=654835 $Y=-7792 $D=0
M1346 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=655525 $Y=-7792 $D=0
M1347 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=656215 $Y=-7792 $D=0
M1348 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=656905 $Y=-7792 $D=0
M1349 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=657595 $Y=-7792 $D=0
M1350 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=658285 $Y=-7792 $D=0
M1351 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=658975 $Y=-7792 $D=0
M1352 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=659665 $Y=-7792 $D=0
M1353 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=660355 $Y=-7792 $D=0
M1354 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=661045 $Y=-7792 $D=0
M1355 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=661735 $Y=-7792 $D=0
M1356 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=662425 $Y=-7792 $D=0
M1357 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=663115 $Y=-7792 $D=0
M1358 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=663805 $Y=-7792 $D=0
M1359 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=664495 $Y=-7792 $D=0
M1360 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=665185 $Y=-7792 $D=0
M1361 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=665875 $Y=-7792 $D=0
M1362 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=666565 $Y=-7792 $D=0
M1363 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=667255 $Y=-7792 $D=0
M1364 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=667945 $Y=-7792 $D=0
M1365 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=668635 $Y=-7792 $D=0
M1366 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=669325 $Y=-7792 $D=0
M1367 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=670015 $Y=-7792 $D=0
M1368 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=670705 $Y=-7792 $D=0
M1369 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=671395 $Y=-7792 $D=0
M1370 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.425e-13 AS=1.275e-13 PD=5.7e-07 PS=5.1e-07 $X=672085 $Y=-7792 $D=0
M1371 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.425e-13 PD=5.1e-07 PS=5.7e-07 $X=672835 $Y=-7792 $D=0
M1372 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=673525 $Y=-7792 $D=0
M1373 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=674215 $Y=-7792 $D=0
M1374 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=674905 $Y=-7792 $D=0
M1375 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=675595 $Y=-7792 $D=0
M1376 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=676285 $Y=-7792 $D=0
M1377 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=676975 $Y=-7792 $D=0
M1378 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=677665 $Y=-7792 $D=0
M1379 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=678355 $Y=-7792 $D=0
M1380 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=679045 $Y=-7792 $D=0
M1381 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=679735 $Y=-7792 $D=0
M1382 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=680425 $Y=-7792 $D=0
M1383 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=681115 $Y=-7792 $D=0
M1384 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=681805 $Y=-7792 $D=0
M1385 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=682495 $Y=-7792 $D=0
M1386 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=683185 $Y=-7792 $D=0
M1387 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=683875 $Y=-7792 $D=0
M1388 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=684565 $Y=-7792 $D=0
M1389 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=685255 $Y=-7792 $D=0
M1390 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=685945 $Y=-7792 $D=0
M1391 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=686635 $Y=-7792 $D=0
M1392 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=687325 $Y=-7792 $D=0
M1393 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=688015 $Y=-7792 $D=0
M1394 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=688705 $Y=-7792 $D=0
M1395 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=689395 $Y=-7792 $D=0
M1396 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=690085 $Y=-7792 $D=0
M1397 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=690775 $Y=-7792 $D=0
M1398 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=691465 $Y=-7792 $D=0
M1399 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=692155 $Y=-7792 $D=0
M1400 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=692845 $Y=-7792 $D=0
M1401 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=693535 $Y=-7792 $D=0
M1402 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=694225 $Y=-7792 $D=0
M1403 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=694915 $Y=-7792 $D=0
M1404 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=695605 $Y=-7792 $D=0
M1405 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=696295 $Y=-7792 $D=0
M1406 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=696985 $Y=-7792 $D=0
M1407 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=697675 $Y=-7792 $D=0
M1408 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=698365 $Y=-7792 $D=0
M1409 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=699055 $Y=-7792 $D=0
M1410 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=699745 $Y=-7792 $D=0
M1411 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=700435 $Y=-7792 $D=0
M1412 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=701125 $Y=-7792 $D=0
M1413 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=701815 $Y=-7792 $D=0
M1414 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=702505 $Y=-7792 $D=0
M1415 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=703195 $Y=-7792 $D=0
M1416 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=703885 $Y=-7792 $D=0
M1417 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=704575 $Y=-7792 $D=0
M1418 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=705265 $Y=-7792 $D=0
M1419 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=705955 $Y=-7792 $D=0
M1420 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=706645 $Y=-7792 $D=0
M1421 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=707335 $Y=-7792 $D=0
M1422 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=708025 $Y=-7792 $D=0
M1423 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=708715 $Y=-7792 $D=0
M1424 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=709405 $Y=-7792 $D=0
M1425 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=710095 $Y=-7792 $D=0
M1426 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=710785 $Y=-7792 $D=0
M1427 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=711475 $Y=-7792 $D=0
M1428 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=712165 $Y=-7792 $D=0
M1429 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=712855 $Y=-7792 $D=0
M1430 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=713545 $Y=-7792 $D=0
M1431 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=714235 $Y=-7792 $D=0
M1432 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=714925 $Y=-7792 $D=0
M1433 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=715615 $Y=-7792 $D=0
M1434 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=716305 $Y=-7792 $D=0
M1435 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=716995 $Y=-7792 $D=0
M1436 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=717685 $Y=-7792 $D=0
M1437 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=718375 $Y=-7792 $D=0
M1438 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=719065 $Y=-7792 $D=0
M1439 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=719755 $Y=-7792 $D=0
M1440 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=720445 $Y=-7792 $D=0
M1441 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=721135 $Y=-7792 $D=0
M1442 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=721825 $Y=-7792 $D=0
M1443 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=722515 $Y=-7792 $D=0
M1444 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=723205 $Y=-7792 $D=0
M1445 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=723895 $Y=-7792 $D=0
M1446 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=724585 $Y=-7792 $D=0
M1447 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=725275 $Y=-7792 $D=0
M1448 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=725965 $Y=-7792 $D=0
M1449 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=726655 $Y=-7792 $D=0
M1450 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=727345 $Y=-7792 $D=0
M1451 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=728035 $Y=-7792 $D=0
M1452 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=728725 $Y=-7792 $D=0
M1453 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=729415 $Y=-7792 $D=0
M1454 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=730105 $Y=-7792 $D=0
M1455 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=730795 $Y=-7792 $D=0
M1456 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=731485 $Y=-7792 $D=0
M1457 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=732175 $Y=-7792 $D=0
M1458 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=732865 $Y=-7792 $D=0
M1459 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=733555 $Y=-7792 $D=0
M1460 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=734245 $Y=-7792 $D=0
M1461 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=734935 $Y=-7792 $D=0
M1462 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=735625 $Y=-7792 $D=0
M1463 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=736315 $Y=-7792 $D=0
M1464 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=737005 $Y=-7792 $D=0
M1465 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=737695 $Y=-7792 $D=0
M1466 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=738385 $Y=-7792 $D=0
M1467 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=739075 $Y=-7792 $D=0
M1468 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=739765 $Y=-7792 $D=0
M1469 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=740455 $Y=-7792 $D=0
M1470 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=741145 $Y=-7792 $D=0
M1471 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=741835 $Y=-7792 $D=0
M1472 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=742525 $Y=-7792 $D=0
M1473 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=743215 $Y=-7792 $D=0
M1474 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=743905 $Y=-7792 $D=0
M1475 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=744595 $Y=-7792 $D=0
M1476 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=745285 $Y=-7792 $D=0
M1477 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=745975 $Y=-7792 $D=0
M1478 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=746665 $Y=-7792 $D=0
M1479 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=747355 $Y=-7792 $D=0
M1480 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=748045 $Y=-7792 $D=0
M1481 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=748735 $Y=-7792 $D=0
M1482 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=749425 $Y=-7792 $D=0
M1483 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=750115 $Y=-7792 $D=0
M1484 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=750805 $Y=-7792 $D=0
M1485 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=751495 $Y=-7792 $D=0
M1486 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=752185 $Y=-7792 $D=0
M1487 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=752875 $Y=-7792 $D=0
M1488 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=753565 $Y=-7792 $D=0
M1489 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=754255 $Y=-7792 $D=0
M1490 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=754945 $Y=-7792 $D=0
M1491 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=755635 $Y=-7792 $D=0
M1492 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=756325 $Y=-7792 $D=0
M1493 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=757015 $Y=-7792 $D=0
M1494 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=757705 $Y=-7792 $D=0
M1495 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=758395 $Y=-7792 $D=0
M1496 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=759085 $Y=-7792 $D=0
M1497 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=759775 $Y=-7792 $D=0
M1498 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=760465 $Y=-7792 $D=0
M1499 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=761155 $Y=-7792 $D=0
M1500 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=761845 $Y=-7792 $D=0
M1501 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=762535 $Y=-7792 $D=0
M1502 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=763225 $Y=-7792 $D=0
M1503 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=763915 $Y=-7792 $D=0
M1504 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=764605 $Y=-7792 $D=0
M1505 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=765295 $Y=-7792 $D=0
M1506 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=765985 $Y=-7792 $D=0
M1507 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=766675 $Y=-7792 $D=0
M1508 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=767365 $Y=-7792 $D=0
M1509 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=768055 $Y=-7792 $D=0
M1510 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=768745 $Y=-7792 $D=0
M1511 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=769435 $Y=-7792 $D=0
M1512 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=770125 $Y=-7792 $D=0
M1513 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=770815 $Y=-7792 $D=0
M1514 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=771505 $Y=-7792 $D=0
M1515 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=772195 $Y=-7792 $D=0
M1516 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=772885 $Y=-7792 $D=0
M1517 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=773575 $Y=-7792 $D=0
M1518 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=774265 $Y=-7792 $D=0
M1519 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=774955 $Y=-7792 $D=0
M1520 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=775645 $Y=-7792 $D=0
M1521 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=776335 $Y=-7792 $D=0
M1522 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=777025 $Y=-7792 $D=0
M1523 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=777715 $Y=-7792 $D=0
M1524 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=778405 $Y=-7792 $D=0
M1525 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=779095 $Y=-7792 $D=0
M1526 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=779785 $Y=-7792 $D=0
M1527 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=780475 $Y=-7792 $D=0
M1528 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=781165 $Y=-7792 $D=0
M1529 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=781855 $Y=-7792 $D=0
M1530 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=782545 $Y=-7792 $D=0
M1531 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=783235 $Y=-7792 $D=0
M1532 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=783925 $Y=-7792 $D=0
M1533 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=784615 $Y=-7792 $D=0
M1534 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=785305 $Y=-7792 $D=0
M1535 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=785995 $Y=-7792 $D=0
M1536 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=786685 $Y=-7792 $D=0
M1537 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=787375 $Y=-7792 $D=0
M1538 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=788065 $Y=-7792 $D=0
M1539 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=788755 $Y=-7792 $D=0
M1540 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=789445 $Y=-7792 $D=0
M1541 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=790135 $Y=-7792 $D=0
M1542 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=790825 $Y=-7792 $D=0
M1543 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=791515 $Y=-7792 $D=0
M1544 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=792205 $Y=-7792 $D=0
M1545 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=792895 $Y=-7792 $D=0
M1546 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=793585 $Y=-7792 $D=0
M1547 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=794275 $Y=-7792 $D=0
M1548 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=794965 $Y=-7792 $D=0
M1549 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=795655 $Y=-7792 $D=0
M1550 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=796345 $Y=-7792 $D=0
M1551 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=797035 $Y=-7792 $D=0
M1552 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=797725 $Y=-7792 $D=0
M1553 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=798415 $Y=-7792 $D=0
M1554 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=799105 $Y=-7792 $D=0
M1555 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=799795 $Y=-7792 $D=0
M1556 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=800485 $Y=-7792 $D=0
M1557 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=801175 $Y=-7792 $D=0
M1558 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=801865 $Y=-7792 $D=0
M1559 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=802555 $Y=-7792 $D=0
M1560 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=803245 $Y=-7792 $D=0
M1561 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=803935 $Y=-7792 $D=0
M1562 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=804625 $Y=-7792 $D=0
M1563 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=805315 $Y=-7792 $D=0
M1564 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=806005 $Y=-7792 $D=0
M1565 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=806695 $Y=-7792 $D=0
M1566 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=807385 $Y=-7792 $D=0
M1567 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=808075 $Y=-7792 $D=0
M1568 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=808765 $Y=-7792 $D=0
M1569 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=809455 $Y=-7792 $D=0
M1570 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=810145 $Y=-7792 $D=0
M1571 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=810835 $Y=-7792 $D=0
M1572 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=811525 $Y=-7792 $D=0
M1573 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=812215 $Y=-7792 $D=0
M1574 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=812905 $Y=-7792 $D=0
M1575 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=813595 $Y=-7792 $D=0
M1576 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=814285 $Y=-7792 $D=0
M1577 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=814975 $Y=-7792 $D=0
M1578 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=815665 $Y=-7792 $D=0
M1579 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=816355 $Y=-7792 $D=0
M1580 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=817045 $Y=-7792 $D=0
M1581 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=817735 $Y=-7792 $D=0
M1582 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=818425 $Y=-7792 $D=0
M1583 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=819115 $Y=-7792 $D=0
M1584 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=819805 $Y=-7792 $D=0
M1585 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=820495 $Y=-7792 $D=0
M1586 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=821185 $Y=-7792 $D=0
M1587 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=821875 $Y=-7792 $D=0
M1588 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=822565 $Y=-7792 $D=0
M1589 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=823255 $Y=-7792 $D=0
M1590 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=823945 $Y=-7792 $D=0
M1591 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=824635 $Y=-7792 $D=0
M1592 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=825325 $Y=-7792 $D=0
M1593 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=826015 $Y=-7792 $D=0
M1594 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=826705 $Y=-7792 $D=0
M1595 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=827395 $Y=-7792 $D=0
M1596 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=828085 $Y=-7792 $D=0
M1597 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=828775 $Y=-7792 $D=0
M1598 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=829465 $Y=-7792 $D=0
M1599 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=830155 $Y=-7792 $D=0
M1600 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=830845 $Y=-7792 $D=0
M1601 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=831535 $Y=-7792 $D=0
M1602 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=832225 $Y=-7792 $D=0
M1603 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=832915 $Y=-7792 $D=0
M1604 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=833605 $Y=-7792 $D=0
M1605 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=834295 $Y=-7792 $D=0
M1606 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=834985 $Y=-7792 $D=0
M1607 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=835675 $Y=-7792 $D=0
M1608 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=836365 $Y=-7792 $D=0
M1609 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=837055 $Y=-7792 $D=0
M1610 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=837745 $Y=-7792 $D=0
M1611 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=838435 $Y=-7792 $D=0
M1612 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=839125 $Y=-7792 $D=0
M1613 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=839815 $Y=-7792 $D=0
M1614 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=840505 $Y=-7792 $D=0
M1615 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=841195 $Y=-7792 $D=0
M1616 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=841885 $Y=-7792 $D=0
M1617 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=842575 $Y=-7792 $D=0
M1618 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=843265 $Y=-7792 $D=0
M1619 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=843955 $Y=-7792 $D=0
M1620 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=844645 $Y=-7792 $D=0
M1621 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=845335 $Y=-7792 $D=0
M1622 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=846025 $Y=-7792 $D=0
M1623 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=846715 $Y=-7792 $D=0
M1624 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=847405 $Y=-7792 $D=0
M1625 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=848095 $Y=-7792 $D=0
M1626 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=848785 $Y=-7792 $D=0
M1627 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=849475 $Y=-7792 $D=0
M1628 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=850165 $Y=-7792 $D=0
M1629 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=850855 $Y=-7792 $D=0
M1630 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=851545 $Y=-7792 $D=0
M1631 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=852235 $Y=-7792 $D=0
M1632 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=852925 $Y=-7792 $D=0
M1633 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=853615 $Y=-7792 $D=0
M1634 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=854305 $Y=-7792 $D=0
M1635 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=854995 $Y=-7792 $D=0
M1636 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=855685 $Y=-7792 $D=0
M1637 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=856375 $Y=-7792 $D=0
M1638 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=857065 $Y=-7792 $D=0
M1639 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=857755 $Y=-7792 $D=0
M1640 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=858445 $Y=-7792 $D=0
M1641 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=859135 $Y=-7792 $D=0
M1642 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=859825 $Y=-7792 $D=0
M1643 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=860515 $Y=-7792 $D=0
M1644 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=861205 $Y=-7792 $D=0
M1645 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=861895 $Y=-7792 $D=0
M1646 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=862585 $Y=-7792 $D=0
M1647 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=863275 $Y=-7792 $D=0
M1648 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=863965 $Y=-7792 $D=0
M1649 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=864655 $Y=-7792 $D=0
M1650 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=865345 $Y=-7792 $D=0
M1651 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=866035 $Y=-7792 $D=0
M1652 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=866725 $Y=-7792 $D=0
M1653 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=867415 $Y=-7792 $D=0
M1654 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=868105 $Y=-7792 $D=0
M1655 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=868795 $Y=-7792 $D=0
M1656 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=869485 $Y=-7792 $D=0
M1657 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=870175 $Y=-7792 $D=0
M1658 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=870865 $Y=-7792 $D=0
M1659 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=871555 $Y=-7792 $D=0
M1660 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=872245 $Y=-7792 $D=0
M1661 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=872935 $Y=-7792 $D=0
M1662 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=873625 $Y=-7792 $D=0
M1663 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=874315 $Y=-7792 $D=0
M1664 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=875005 $Y=-7792 $D=0
M1665 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=875695 $Y=-7792 $D=0
M1666 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=876385 $Y=-7792 $D=0
M1667 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=877075 $Y=-7792 $D=0
M1668 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=877765 $Y=-7792 $D=0
M1669 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=878455 $Y=-7792 $D=0
M1670 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=879145 $Y=-7792 $D=0
M1671 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=879835 $Y=-7792 $D=0
M1672 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=880525 $Y=-7792 $D=0
M1673 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=881215 $Y=-7792 $D=0
M1674 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=881905 $Y=-7792 $D=0
M1675 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=882595 $Y=-7792 $D=0
M1676 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=883285 $Y=-7792 $D=0
M1677 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=883975 $Y=-7792 $D=0
M1678 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=884665 $Y=-7792 $D=0
M1679 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=885355 $Y=-7792 $D=0
M1680 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=886045 $Y=-7792 $D=0
M1681 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=886735 $Y=-7792 $D=0
M1682 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=887425 $Y=-7792 $D=0
M1683 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=888115 $Y=-7792 $D=0
M1684 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=888805 $Y=-7792 $D=0
M1685 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=889495 $Y=-7792 $D=0
M1686 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=890185 $Y=-7792 $D=0
M1687 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=890875 $Y=-7792 $D=0
M1688 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=891565 $Y=-7792 $D=0
M1689 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=892255 $Y=-7792 $D=0
M1690 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=892945 $Y=-7792 $D=0
M1691 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=893635 $Y=-7792 $D=0
M1692 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=894325 $Y=-7792 $D=0
M1693 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=895015 $Y=-7792 $D=0
M1694 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=895705 $Y=-7792 $D=0
M1695 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=896395 $Y=-7792 $D=0
M1696 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=897085 $Y=-7792 $D=0
M1697 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=897775 $Y=-7792 $D=0
M1698 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=898465 $Y=-7792 $D=0
M1699 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=899155 $Y=-7792 $D=0
M1700 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=899845 $Y=-7792 $D=0
M1701 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=900535 $Y=-7792 $D=0
M1702 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=901225 $Y=-7792 $D=0
M1703 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=901915 $Y=-7792 $D=0
M1704 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=902605 $Y=-7792 $D=0
M1705 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=903295 $Y=-7792 $D=0
M1706 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=903985 $Y=-7792 $D=0
M1707 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=904675 $Y=-7792 $D=0
M1708 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=905365 $Y=-7792 $D=0
M1709 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=906055 $Y=-7792 $D=0
M1710 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=906745 $Y=-7792 $D=0
M1711 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=907435 $Y=-7792 $D=0
M1712 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=908125 $Y=-7792 $D=0
M1713 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=908815 $Y=-7792 $D=0
M1714 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=909505 $Y=-7792 $D=0
M1715 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=910195 $Y=-7792 $D=0
M1716 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=910885 $Y=-7792 $D=0
M1717 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=911575 $Y=-7792 $D=0
M1718 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=912265 $Y=-7792 $D=0
M1719 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=912955 $Y=-7792 $D=0
M1720 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=913645 $Y=-7792 $D=0
M1721 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=914335 $Y=-7792 $D=0
M1722 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=915025 $Y=-7792 $D=0
M1723 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=915715 $Y=-7792 $D=0
M1724 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=916405 $Y=-7792 $D=0
M1725 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=917095 $Y=-7792 $D=0
M1726 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=917785 $Y=-7792 $D=0
M1727 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=918475 $Y=-7792 $D=0
M1728 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=919165 $Y=-7792 $D=0
M1729 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=919855 $Y=-7792 $D=0
M1730 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=920545 $Y=-7792 $D=0
M1731 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=921235 $Y=-7792 $D=0
M1732 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=921925 $Y=-7792 $D=0
M1733 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=922615 $Y=-7792 $D=0
M1734 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=923305 $Y=-7792 $D=0
M1735 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=923995 $Y=-7792 $D=0
M1736 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=924685 $Y=-7792 $D=0
M1737 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=925375 $Y=-7792 $D=0
M1738 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=926065 $Y=-7792 $D=0
M1739 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=926755 $Y=-7792 $D=0
M1740 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=927445 $Y=-7792 $D=0
M1741 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=928135 $Y=-7792 $D=0
M1742 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=928825 $Y=-7792 $D=0
M1743 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=929515 $Y=-7792 $D=0
M1744 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=930205 $Y=-7792 $D=0
M1745 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=930895 $Y=-7792 $D=0
M1746 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=931585 $Y=-7792 $D=0
M1747 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=932275 $Y=-7792 $D=0
M1748 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=932965 $Y=-7792 $D=0
M1749 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=933655 $Y=-7792 $D=0
M1750 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=934345 $Y=-7792 $D=0
M1751 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=935035 $Y=-7792 $D=0
M1752 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=935725 $Y=-7792 $D=0
M1753 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=936415 $Y=-7792 $D=0
M1754 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=937105 $Y=-7792 $D=0
M1755 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=937795 $Y=-7792 $D=0
M1756 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=938485 $Y=-7792 $D=0
M1757 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=939175 $Y=-7792 $D=0
M1758 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=939865 $Y=-7792 $D=0
M1759 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=940555 $Y=-7792 $D=0
M1760 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=941245 $Y=-7792 $D=0
M1761 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=941935 $Y=-7792 $D=0
M1762 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=942625 $Y=-7792 $D=0
M1763 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=943315 $Y=-7792 $D=0
M1764 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=944005 $Y=-7792 $D=0
M1765 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=944695 $Y=-7792 $D=0
M1766 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=945385 $Y=-7792 $D=0
M1767 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=946075 $Y=-7792 $D=0
M1768 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=946765 $Y=-7792 $D=0
M1769 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=947455 $Y=-7792 $D=0
M1770 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=948145 $Y=-7792 $D=0
M1771 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=948835 $Y=-7792 $D=0
M1772 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=949525 $Y=-7792 $D=0
M1773 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=950215 $Y=-7792 $D=0
M1774 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=950905 $Y=-7792 $D=0
M1775 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=951595 $Y=-7792 $D=0
M1776 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=952285 $Y=-7792 $D=0
M1777 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=952975 $Y=-7792 $D=0
M1778 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=953665 $Y=-7792 $D=0
M1779 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=954355 $Y=-7792 $D=0
M1780 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=955045 $Y=-7792 $D=0
M1781 Vcout 19 GND GND N_18 L=1.8e-07 W=5e-07 AD=1.275e-13 AS=1.275e-13 PD=5.1e-07 PS=5.1e-07 $X=955735 $Y=-7792 $D=0
M1782 GND 19 Vcout GND N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.275e-13 PD=1.48e-06 PS=5.1e-07 $X=956425 $Y=-7792 $D=0
M1783 4 Vin VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=9.0454e-13 PD=2.826e-06 PS=2.826e-06 $X=-145 $Y=1334 $D=1
M1784 5 4 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=1415 $Y=1334 $D=1
M1785 VDD 4 5 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=2105 $Y=1334 $D=1
M1786 5 4 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=2795 $Y=1334 $D=1
M1787 VDD 4 5 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=3485 $Y=1334 $D=1
M1788 5 4 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=4175 $Y=1334 $D=1
M1789 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=5735 $Y=1334 $D=1
M1790 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=6425 $Y=1334 $D=1
M1791 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=7115 $Y=1334 $D=1
M1792 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=7805 $Y=1334 $D=1
M1793 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=8495 $Y=1334 $D=1
M1794 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=9185 $Y=1334 $D=1
M1795 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=9875 $Y=1334 $D=1
M1796 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=10565 $Y=1334 $D=1
M1797 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=11255 $Y=1334 $D=1
M1798 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=11945 $Y=1334 $D=1
M1799 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=12635 $Y=1334 $D=1
M1800 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=13325 $Y=1334 $D=1
M1801 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=14015 $Y=1334 $D=1
M1802 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=14705 $Y=1334 $D=1
M1803 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=15395 $Y=1334 $D=1
M1804 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=16085 $Y=1334 $D=1
M1805 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=16775 $Y=1334 $D=1
M1806 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=17465 $Y=1334 $D=1
M1807 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=18155 $Y=1334 $D=1
M1808 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=18845 $Y=1334 $D=1
M1809 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=19535 $Y=1334 $D=1
M1810 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=20225 $Y=1334 $D=1
M1811 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=20915 $Y=1334 $D=1
M1812 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=21605 $Y=1334 $D=1
M1813 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=22295 $Y=1334 $D=1
M1814 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=22985 $Y=1334 $D=1
M1815 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=23675 $Y=1334 $D=1
M1816 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=24365 $Y=1334 $D=1
M1817 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=25055 $Y=1334 $D=1
M1818 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=25745 $Y=1334 $D=1
M1819 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=26435 $Y=1334 $D=1
M1820 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=27125 $Y=1334 $D=1
M1821 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=27815 $Y=1334 $D=1
M1822 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=28505 $Y=1334 $D=1
M1823 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=29195 $Y=1334 $D=1
M1824 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=29885 $Y=1334 $D=1
M1825 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=30575 $Y=1334 $D=1
M1826 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=31265 $Y=1334 $D=1
M1827 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=31955 $Y=1334 $D=1
M1828 VDD 5 6 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=32645 $Y=1334 $D=1
M1829 6 5 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=33335 $Y=1334 $D=1
M1830 7 6 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=9.0454e-13 PD=2.826e-06 PS=2.826e-06 $X=38665 $Y=-6292 $D=1
M1831 8 6 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=9.0454e-13 PD=2.826e-06 PS=2.826e-06 $X=38665 $Y=1334 $D=1
M1832 9 6 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=9.0454e-13 PD=2.826e-06 PS=2.826e-06 $X=38665 $Y=8960 $D=1
M1833 10 7 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=40225 $Y=-6292 $D=1
M1834 11 8 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=40225 $Y=1334 $D=1
M1835 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=40225 $Y=8960 $D=1
M1836 VDD 7 10 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=40915 $Y=-6292 $D=1
M1837 VDD 8 11 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=40915 $Y=1334 $D=1
M1838 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=40915 $Y=8960 $D=1
M1839 10 7 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=41605 $Y=-6292 $D=1
M1840 11 8 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=41605 $Y=1334 $D=1
M1841 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=41605 $Y=8960 $D=1
M1842 VDD 8 11 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=42295 $Y=1334 $D=1
M1843 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=42295 $Y=8960 $D=1
M1844 11 8 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=42985 $Y=1334 $D=1
M1845 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=42985 $Y=8960 $D=1
M1846 12 10 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=43165 $Y=-6292 $D=1
M1847 VDD 8 11 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=43675 $Y=1334 $D=1
M1848 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=43675 $Y=8960 $D=1
M1849 VDD 10 12 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=43855 $Y=-6292 $D=1
M1850 11 8 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=44365 $Y=1334 $D=1
M1851 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=44365 $Y=8960 $D=1
M1852 12 10 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=44545 $Y=-6292 $D=1
M1853 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=45055 $Y=8960 $D=1
M1854 VDD 10 12 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=45235 $Y=-6292 $D=1
M1855 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=45745 $Y=8960 $D=1
M1856 12 10 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=45925 $Y=-6292 $D=1
M1857 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=45925 $Y=1334 $D=1
M1858 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=46435 $Y=8960 $D=1
M1859 VDD 10 12 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=46615 $Y=-6292 $D=1
M1860 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=46615 $Y=1334 $D=1
M1861 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=47125 $Y=8960 $D=1
M1862 12 10 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=47305 $Y=-6292 $D=1
M1863 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=47305 $Y=1334 $D=1
M1864 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=47815 $Y=8960 $D=1
M1865 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=47995 $Y=1334 $D=1
M1866 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=48505 $Y=8960 $D=1
M1867 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=48685 $Y=1334 $D=1
M1868 13 12 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=48865 $Y=-6292 $D=1
M1869 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=49195 $Y=8960 $D=1
M1870 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=49375 $Y=1334 $D=1
M1871 VDD 12 13 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=49555 $Y=-6292 $D=1
M1872 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=49885 $Y=8960 $D=1
M1873 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=50065 $Y=1334 $D=1
M1874 13 12 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=50245 $Y=-6292 $D=1
M1875 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=50575 $Y=8960 $D=1
M1876 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=50755 $Y=1334 $D=1
M1877 VDD 12 13 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=50935 $Y=-6292 $D=1
M1878 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=51265 $Y=8960 $D=1
M1879 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=51445 $Y=1334 $D=1
M1880 13 12 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=51625 $Y=-6292 $D=1
M1881 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=51955 $Y=8960 $D=1
M1882 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=52135 $Y=1334 $D=1
M1883 VDD 12 13 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=52315 $Y=-6292 $D=1
M1884 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=52645 $Y=8960 $D=1
M1885 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=52825 $Y=1334 $D=1
M1886 13 12 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=53005 $Y=-6292 $D=1
M1887 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=53335 $Y=8960 $D=1
M1888 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=53515 $Y=1334 $D=1
M1889 VDD 12 13 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=53695 $Y=-6292 $D=1
M1890 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=54025 $Y=8960 $D=1
M1891 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=54205 $Y=1334 $D=1
M1892 13 12 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=54385 $Y=-6292 $D=1
M1893 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=54715 $Y=8960 $D=1
M1894 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=54895 $Y=1334 $D=1
M1895 VDD 12 13 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=55075 $Y=-6292 $D=1
M1896 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=55405 $Y=8960 $D=1
M1897 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=55585 $Y=1334 $D=1
M1898 13 12 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=55765 $Y=-6292 $D=1
M1899 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=56095 $Y=8960 $D=1
M1900 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=56275 $Y=1334 $D=1
M1901 VDD 12 13 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=56455 $Y=-6292 $D=1
M1902 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=56785 $Y=8960 $D=1
M1903 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=56965 $Y=1334 $D=1
M1904 13 12 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=57145 $Y=-6292 $D=1
M1905 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=57475 $Y=8960 $D=1
M1906 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=57655 $Y=1334 $D=1
M1907 VDD 12 13 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=57835 $Y=-6292 $D=1
M1908 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=58165 $Y=8960 $D=1
M1909 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=58345 $Y=1334 $D=1
M1910 13 12 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=58525 $Y=-6292 $D=1
M1911 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=58855 $Y=8960 $D=1
M1912 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=59035 $Y=1334 $D=1
M1913 VDD 12 13 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=59215 $Y=-6292 $D=1
M1914 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=59545 $Y=8960 $D=1
M1915 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=59725 $Y=1334 $D=1
M1916 13 12 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=59905 $Y=-6292 $D=1
M1917 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=60235 $Y=8960 $D=1
M1918 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=60415 $Y=1334 $D=1
M1919 VDD 12 13 VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=60595 $Y=-6292 $D=1
M1920 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=60925 $Y=8960 $D=1
M1921 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=61105 $Y=1334 $D=1
M1922 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=61615 $Y=8960 $D=1
M1923 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=61795 $Y=1334 $D=1
M1924 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=62155 $Y=-6292 $D=1
M1925 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=62305 $Y=8960 $D=1
M1926 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=62485 $Y=1334 $D=1
M1927 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=62845 $Y=-6292 $D=1
M1928 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=62995 $Y=8960 $D=1
M1929 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=63175 $Y=1334 $D=1
M1930 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=63535 $Y=-6292 $D=1
M1931 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=63685 $Y=8960 $D=1
M1932 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=63865 $Y=1334 $D=1
M1933 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=64225 $Y=-6292 $D=1
M1934 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=64375 $Y=8960 $D=1
M1935 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=64555 $Y=1334 $D=1
M1936 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=64915 $Y=-6292 $D=1
M1937 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=65065 $Y=8960 $D=1
M1938 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=65245 $Y=1334 $D=1
M1939 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=65605 $Y=-6292 $D=1
M1940 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=65755 $Y=8960 $D=1
M1941 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=65935 $Y=1334 $D=1
M1942 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=66295 $Y=-6292 $D=1
M1943 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=66445 $Y=8960 $D=1
M1944 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=66625 $Y=1334 $D=1
M1945 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=66985 $Y=-6292 $D=1
M1946 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=67135 $Y=8960 $D=1
M1947 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=67315 $Y=1334 $D=1
M1948 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=67675 $Y=-6292 $D=1
M1949 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=67825 $Y=8960 $D=1
M1950 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=68005 $Y=1334 $D=1
M1951 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=68365 $Y=-6292 $D=1
M1952 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=68515 $Y=8960 $D=1
M1953 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=68695 $Y=1334 $D=1
M1954 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=69055 $Y=-6292 $D=1
M1955 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=69205 $Y=8960 $D=1
M1956 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=69385 $Y=1334 $D=1
M1957 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=69745 $Y=-6292 $D=1
M1958 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=69895 $Y=8960 $D=1
M1959 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=70075 $Y=1334 $D=1
M1960 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=70435 $Y=-6292 $D=1
M1961 Vaout 9 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=70585 $Y=8960 $D=1
M1962 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=70765 $Y=1334 $D=1
M1963 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=71125 $Y=-6292 $D=1
M1964 VDD 9 Vaout VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=71275 $Y=8960 $D=1
M1965 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=71455 $Y=1334 $D=1
M1966 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=71815 $Y=-6292 $D=1
M1967 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=72145 $Y=1334 $D=1
M1968 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=72505 $Y=-6292 $D=1
M1969 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=72835 $Y=1334 $D=1
M1970 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=73195 $Y=-6292 $D=1
M1971 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=73525 $Y=1334 $D=1
M1972 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=73885 $Y=-6292 $D=1
M1973 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=74215 $Y=1334 $D=1
M1974 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=74575 $Y=-6292 $D=1
M1975 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=74905 $Y=1334 $D=1
M1976 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=75265 $Y=-6292 $D=1
M1977 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=75595 $Y=1334 $D=1
M1978 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=75955 $Y=-6292 $D=1
M1979 15 11 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=76285 $Y=1334 $D=1
M1980 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=76645 $Y=-6292 $D=1
M1981 VDD 11 15 VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=76975 $Y=1334 $D=1
M1982 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=77335 $Y=-6292 $D=1
M1983 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=78025 $Y=-6292 $D=1
M1984 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=78535 $Y=1334 $D=1
M1985 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=78715 $Y=-6292 $D=1
M1986 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=79225 $Y=1334 $D=1
M1987 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=79405 $Y=-6292 $D=1
M1988 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=79915 $Y=1334 $D=1
M1989 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=80095 $Y=-6292 $D=1
M1990 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=80605 $Y=1334 $D=1
M1991 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=80785 $Y=-6292 $D=1
M1992 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=81295 $Y=1334 $D=1
M1993 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=81475 $Y=-6292 $D=1
M1994 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=81985 $Y=1334 $D=1
M1995 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=82165 $Y=-6292 $D=1
M1996 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=82675 $Y=1334 $D=1
M1997 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=82855 $Y=-6292 $D=1
M1998 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=83365 $Y=1334 $D=1
M1999 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=83545 $Y=-6292 $D=1
M2000 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=84055 $Y=1334 $D=1
M2001 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=84235 $Y=-6292 $D=1
M2002 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=84745 $Y=1334 $D=1
M2003 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=84925 $Y=-6292 $D=1
M2004 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=85435 $Y=1334 $D=1
M2005 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=85615 $Y=-6292 $D=1
M2006 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=86125 $Y=1334 $D=1
M2007 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=86305 $Y=-6292 $D=1
M2008 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=86815 $Y=1334 $D=1
M2009 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=86995 $Y=-6292 $D=1
M2010 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=87505 $Y=1334 $D=1
M2011 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=87685 $Y=-6292 $D=1
M2012 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=88195 $Y=1334 $D=1
M2013 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=88375 $Y=-6292 $D=1
M2014 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=88885 $Y=1334 $D=1
M2015 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=89065 $Y=-6292 $D=1
M2016 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=89575 $Y=1334 $D=1
M2017 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=89755 $Y=-6292 $D=1
M2018 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=90265 $Y=1334 $D=1
M2019 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=90445 $Y=-6292 $D=1
M2020 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=90955 $Y=1334 $D=1
M2021 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=91135 $Y=-6292 $D=1
M2022 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=91645 $Y=1334 $D=1
M2023 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=91825 $Y=-6292 $D=1
M2024 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=92335 $Y=1334 $D=1
M2025 16 13 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=92515 $Y=-6292 $D=1
M2026 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=93025 $Y=1334 $D=1
M2027 VDD 13 16 VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=93205 $Y=-6292 $D=1
M2028 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=93715 $Y=1334 $D=1
M2029 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=94405 $Y=1334 $D=1
M2030 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=94765 $Y=-6292 $D=1
M2031 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=95095 $Y=1334 $D=1
M2032 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=95455 $Y=-6292 $D=1
M2033 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=95785 $Y=1334 $D=1
M2034 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=96145 $Y=-6292 $D=1
M2035 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=96475 $Y=1334 $D=1
M2036 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=96835 $Y=-6292 $D=1
M2037 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=97165 $Y=1334 $D=1
M2038 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=97525 $Y=-6292 $D=1
M2039 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=97855 $Y=1334 $D=1
M2040 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=98215 $Y=-6292 $D=1
M2041 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=98545 $Y=1334 $D=1
M2042 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=98905 $Y=-6292 $D=1
M2043 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=99235 $Y=1334 $D=1
M2044 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=99595 $Y=-6292 $D=1
M2045 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=99925 $Y=1334 $D=1
M2046 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=100285 $Y=-6292 $D=1
M2047 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=100615 $Y=1334 $D=1
M2048 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=100975 $Y=-6292 $D=1
M2049 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=101305 $Y=1334 $D=1
M2050 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=101665 $Y=-6292 $D=1
M2051 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=101995 $Y=1334 $D=1
M2052 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=102355 $Y=-6292 $D=1
M2053 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=102685 $Y=1334 $D=1
M2054 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=103045 $Y=-6292 $D=1
M2055 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=103375 $Y=1334 $D=1
M2056 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=103735 $Y=-6292 $D=1
M2057 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=104065 $Y=1334 $D=1
M2058 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=104425 $Y=-6292 $D=1
M2059 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=104755 $Y=1334 $D=1
M2060 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=105115 $Y=-6292 $D=1
M2061 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=105445 $Y=1334 $D=1
M2062 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=105805 $Y=-6292 $D=1
M2063 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=106135 $Y=1334 $D=1
M2064 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=106495 $Y=-6292 $D=1
M2065 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=106825 $Y=1334 $D=1
M2066 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=107185 $Y=-6292 $D=1
M2067 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=107515 $Y=1334 $D=1
M2068 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=107875 $Y=-6292 $D=1
M2069 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=108205 $Y=1334 $D=1
M2070 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=108565 $Y=-6292 $D=1
M2071 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=108895 $Y=1334 $D=1
M2072 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=109255 $Y=-6292 $D=1
M2073 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=109585 $Y=1334 $D=1
M2074 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=109945 $Y=-6292 $D=1
M2075 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=110275 $Y=1334 $D=1
M2076 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=110635 $Y=-6292 $D=1
M2077 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=110965 $Y=1334 $D=1
M2078 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=111325 $Y=-6292 $D=1
M2079 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=111655 $Y=1334 $D=1
M2080 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=112015 $Y=-6292 $D=1
M2081 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=112345 $Y=1334 $D=1
M2082 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=112705 $Y=-6292 $D=1
M2083 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=113035 $Y=1334 $D=1
M2084 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=113395 $Y=-6292 $D=1
M2085 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=113725 $Y=1334 $D=1
M2086 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=114085 $Y=-6292 $D=1
M2087 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=114415 $Y=1334 $D=1
M2088 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=114775 $Y=-6292 $D=1
M2089 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=115105 $Y=1334 $D=1
M2090 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=115465 $Y=-6292 $D=1
M2091 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=115795 $Y=1334 $D=1
M2092 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=116155 $Y=-6292 $D=1
M2093 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=116485 $Y=1334 $D=1
M2094 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=116845 $Y=-6292 $D=1
M2095 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=117175 $Y=1334 $D=1
M2096 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=117535 $Y=-6292 $D=1
M2097 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=117865 $Y=1334 $D=1
M2098 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=118225 $Y=-6292 $D=1
M2099 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=118555 $Y=1334 $D=1
M2100 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=118915 $Y=-6292 $D=1
M2101 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=119245 $Y=1334 $D=1
M2102 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=119605 $Y=-6292 $D=1
M2103 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=119935 $Y=1334 $D=1
M2104 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=120295 $Y=-6292 $D=1
M2105 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=120625 $Y=1334 $D=1
M2106 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=120985 $Y=-6292 $D=1
M2107 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=121315 $Y=1334 $D=1
M2108 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=121675 $Y=-6292 $D=1
M2109 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=122005 $Y=1334 $D=1
M2110 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=122365 $Y=-6292 $D=1
M2111 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=122695 $Y=1334 $D=1
M2112 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=123055 $Y=-6292 $D=1
M2113 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=123385 $Y=1334 $D=1
M2114 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=123745 $Y=-6292 $D=1
M2115 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=124075 $Y=1334 $D=1
M2116 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=124435 $Y=-6292 $D=1
M2117 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=124765 $Y=1334 $D=1
M2118 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=125125 $Y=-6292 $D=1
M2119 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=125455 $Y=1334 $D=1
M2120 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=125815 $Y=-6292 $D=1
M2121 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=126145 $Y=1334 $D=1
M2122 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=126505 $Y=-6292 $D=1
M2123 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=126835 $Y=1334 $D=1
M2124 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=127195 $Y=-6292 $D=1
M2125 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=127525 $Y=1334 $D=1
M2126 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=127885 $Y=-6292 $D=1
M2127 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=128215 $Y=1334 $D=1
M2128 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=128575 $Y=-6292 $D=1
M2129 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=128905 $Y=1334 $D=1
M2130 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=129265 $Y=-6292 $D=1
M2131 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=129595 $Y=1334 $D=1
M2132 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=129955 $Y=-6292 $D=1
M2133 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=130285 $Y=1334 $D=1
M2134 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=130645 $Y=-6292 $D=1
M2135 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=130975 $Y=1334 $D=1
M2136 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=131335 $Y=-6292 $D=1
M2137 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=131665 $Y=1334 $D=1
M2138 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=132025 $Y=-6292 $D=1
M2139 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=132355 $Y=1334 $D=1
M2140 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=132715 $Y=-6292 $D=1
M2141 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=133045 $Y=1334 $D=1
M2142 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=133405 $Y=-6292 $D=1
M2143 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=133735 $Y=1334 $D=1
M2144 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=134095 $Y=-6292 $D=1
M2145 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=134425 $Y=1334 $D=1
M2146 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=134785 $Y=-6292 $D=1
M2147 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=135115 $Y=1334 $D=1
M2148 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=135475 $Y=-6292 $D=1
M2149 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=135805 $Y=1334 $D=1
M2150 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=136165 $Y=-6292 $D=1
M2151 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=136495 $Y=1334 $D=1
M2152 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=136855 $Y=-6292 $D=1
M2153 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=137185 $Y=1334 $D=1
M2154 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=137545 $Y=-6292 $D=1
M2155 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=137875 $Y=1334 $D=1
M2156 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=138235 $Y=-6292 $D=1
M2157 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=138565 $Y=1334 $D=1
M2158 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=138925 $Y=-6292 $D=1
M2159 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=139255 $Y=1334 $D=1
M2160 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=139615 $Y=-6292 $D=1
M2161 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=5.2611e-13 AS=4.7073e-13 PD=5.7e-07 PS=5.1e-07 $X=139945 $Y=1334 $D=1
M2162 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=140305 $Y=-6292 $D=1
M2163 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=5.2611e-13 PD=5.1e-07 PS=5.7e-07 $X=140695 $Y=1334 $D=1
M2164 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=140995 $Y=-6292 $D=1
M2165 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=141385 $Y=1334 $D=1
M2166 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=141685 $Y=-6292 $D=1
M2167 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=142075 $Y=1334 $D=1
M2168 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=142375 $Y=-6292 $D=1
M2169 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=142765 $Y=1334 $D=1
M2170 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=143065 $Y=-6292 $D=1
M2171 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=143455 $Y=1334 $D=1
M2172 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=143755 $Y=-6292 $D=1
M2173 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=144145 $Y=1334 $D=1
M2174 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=144445 $Y=-6292 $D=1
M2175 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=144835 $Y=1334 $D=1
M2176 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=145135 $Y=-6292 $D=1
M2177 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=145525 $Y=1334 $D=1
M2178 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=145825 $Y=-6292 $D=1
M2179 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=146215 $Y=1334 $D=1
M2180 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=146515 $Y=-6292 $D=1
M2181 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=146905 $Y=1334 $D=1
M2182 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=147205 $Y=-6292 $D=1
M2183 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=147595 $Y=1334 $D=1
M2184 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=147895 $Y=-6292 $D=1
M2185 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=148285 $Y=1334 $D=1
M2186 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=148585 $Y=-6292 $D=1
M2187 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=148975 $Y=1334 $D=1
M2188 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=149275 $Y=-6292 $D=1
M2189 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=149665 $Y=1334 $D=1
M2190 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=149965 $Y=-6292 $D=1
M2191 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=150355 $Y=1334 $D=1
M2192 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=150655 $Y=-6292 $D=1
M2193 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=151045 $Y=1334 $D=1
M2194 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=151345 $Y=-6292 $D=1
M2195 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=151735 $Y=1334 $D=1
M2196 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=152035 $Y=-6292 $D=1
M2197 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=152425 $Y=1334 $D=1
M2198 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=152725 $Y=-6292 $D=1
M2199 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=153115 $Y=1334 $D=1
M2200 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=153415 $Y=-6292 $D=1
M2201 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=153805 $Y=1334 $D=1
M2202 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=154105 $Y=-6292 $D=1
M2203 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=154495 $Y=1334 $D=1
M2204 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=154795 $Y=-6292 $D=1
M2205 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=155185 $Y=1334 $D=1
M2206 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=155485 $Y=-6292 $D=1
M2207 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=155875 $Y=1334 $D=1
M2208 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=156175 $Y=-6292 $D=1
M2209 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=156565 $Y=1334 $D=1
M2210 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=156865 $Y=-6292 $D=1
M2211 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=157255 $Y=1334 $D=1
M2212 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=157555 $Y=-6292 $D=1
M2213 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=157945 $Y=1334 $D=1
M2214 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=158245 $Y=-6292 $D=1
M2215 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=158635 $Y=1334 $D=1
M2216 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=158935 $Y=-6292 $D=1
M2217 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=159325 $Y=1334 $D=1
M2218 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=159625 $Y=-6292 $D=1
M2219 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=160015 $Y=1334 $D=1
M2220 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=160315 $Y=-6292 $D=1
M2221 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=160705 $Y=1334 $D=1
M2222 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=161005 $Y=-6292 $D=1
M2223 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=161395 $Y=1334 $D=1
M2224 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=161695 $Y=-6292 $D=1
M2225 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=162085 $Y=1334 $D=1
M2226 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=162385 $Y=-6292 $D=1
M2227 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=162775 $Y=1334 $D=1
M2228 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=163075 $Y=-6292 $D=1
M2229 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=163465 $Y=1334 $D=1
M2230 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=163765 $Y=-6292 $D=1
M2231 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=164155 $Y=1334 $D=1
M2232 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=164455 $Y=-6292 $D=1
M2233 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=164845 $Y=1334 $D=1
M2234 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=165145 $Y=-6292 $D=1
M2235 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=165535 $Y=1334 $D=1
M2236 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=165835 $Y=-6292 $D=1
M2237 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=166225 $Y=1334 $D=1
M2238 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=166525 $Y=-6292 $D=1
M2239 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=166915 $Y=1334 $D=1
M2240 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=167215 $Y=-6292 $D=1
M2241 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=167605 $Y=1334 $D=1
M2242 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=167905 $Y=-6292 $D=1
M2243 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=168295 $Y=1334 $D=1
M2244 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=168595 $Y=-6292 $D=1
M2245 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=168985 $Y=1334 $D=1
M2246 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=169285 $Y=-6292 $D=1
M2247 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=169675 $Y=1334 $D=1
M2248 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=169975 $Y=-6292 $D=1
M2249 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=170365 $Y=1334 $D=1
M2250 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=170665 $Y=-6292 $D=1
M2251 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=171055 $Y=1334 $D=1
M2252 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=171355 $Y=-6292 $D=1
M2253 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=171745 $Y=1334 $D=1
M2254 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=172045 $Y=-6292 $D=1
M2255 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=172435 $Y=1334 $D=1
M2256 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=172735 $Y=-6292 $D=1
M2257 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=173125 $Y=1334 $D=1
M2258 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=173425 $Y=-6292 $D=1
M2259 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=173815 $Y=1334 $D=1
M2260 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=174115 $Y=-6292 $D=1
M2261 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=174505 $Y=1334 $D=1
M2262 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=174805 $Y=-6292 $D=1
M2263 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=175195 $Y=1334 $D=1
M2264 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=175495 $Y=-6292 $D=1
M2265 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=175885 $Y=1334 $D=1
M2266 17 16 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=176185 $Y=-6292 $D=1
M2267 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=176575 $Y=1334 $D=1
M2268 VDD 16 17 VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=176875 $Y=-6292 $D=1
M2269 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=177265 $Y=1334 $D=1
M2270 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=177955 $Y=1334 $D=1
M2271 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=178435 $Y=-6292 $D=1
M2272 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=178645 $Y=1334 $D=1
M2273 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=179125 $Y=-6292 $D=1
M2274 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=179335 $Y=1334 $D=1
M2275 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=179815 $Y=-6292 $D=1
M2276 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=180025 $Y=1334 $D=1
M2277 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=180505 $Y=-6292 $D=1
M2278 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=180715 $Y=1334 $D=1
M2279 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=181195 $Y=-6292 $D=1
M2280 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=181405 $Y=1334 $D=1
M2281 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=181885 $Y=-6292 $D=1
M2282 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=182095 $Y=1334 $D=1
M2283 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=182575 $Y=-6292 $D=1
M2284 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=182785 $Y=1334 $D=1
M2285 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=183265 $Y=-6292 $D=1
M2286 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=183475 $Y=1334 $D=1
M2287 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=183955 $Y=-6292 $D=1
M2288 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=184165 $Y=1334 $D=1
M2289 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=184645 $Y=-6292 $D=1
M2290 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=184855 $Y=1334 $D=1
M2291 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=185335 $Y=-6292 $D=1
M2292 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=185545 $Y=1334 $D=1
M2293 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=186025 $Y=-6292 $D=1
M2294 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=186235 $Y=1334 $D=1
M2295 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=186715 $Y=-6292 $D=1
M2296 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=186925 $Y=1334 $D=1
M2297 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=187405 $Y=-6292 $D=1
M2298 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=187615 $Y=1334 $D=1
M2299 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=188095 $Y=-6292 $D=1
M2300 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=188305 $Y=1334 $D=1
M2301 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=188785 $Y=-6292 $D=1
M2302 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=188995 $Y=1334 $D=1
M2303 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=189475 $Y=-6292 $D=1
M2304 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=189685 $Y=1334 $D=1
M2305 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=190165 $Y=-6292 $D=1
M2306 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=190375 $Y=1334 $D=1
M2307 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=190855 $Y=-6292 $D=1
M2308 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=191065 $Y=1334 $D=1
M2309 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=191545 $Y=-6292 $D=1
M2310 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=191755 $Y=1334 $D=1
M2311 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=192235 $Y=-6292 $D=1
M2312 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=192445 $Y=1334 $D=1
M2313 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=192925 $Y=-6292 $D=1
M2314 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=193135 $Y=1334 $D=1
M2315 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=193615 $Y=-6292 $D=1
M2316 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=193825 $Y=1334 $D=1
M2317 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=194305 $Y=-6292 $D=1
M2318 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=194515 $Y=1334 $D=1
M2319 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=194995 $Y=-6292 $D=1
M2320 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=195205 $Y=1334 $D=1
M2321 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=195685 $Y=-6292 $D=1
M2322 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=195895 $Y=1334 $D=1
M2323 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=196375 $Y=-6292 $D=1
M2324 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=196585 $Y=1334 $D=1
M2325 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=197065 $Y=-6292 $D=1
M2326 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=197275 $Y=1334 $D=1
M2327 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=197755 $Y=-6292 $D=1
M2328 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=197965 $Y=1334 $D=1
M2329 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=198445 $Y=-6292 $D=1
M2330 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=198655 $Y=1334 $D=1
M2331 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=199135 $Y=-6292 $D=1
M2332 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=199345 $Y=1334 $D=1
M2333 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=199825 $Y=-6292 $D=1
M2334 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=200035 $Y=1334 $D=1
M2335 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=200515 $Y=-6292 $D=1
M2336 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=200725 $Y=1334 $D=1
M2337 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=201205 $Y=-6292 $D=1
M2338 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=201415 $Y=1334 $D=1
M2339 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=201895 $Y=-6292 $D=1
M2340 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=202105 $Y=1334 $D=1
M2341 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=202585 $Y=-6292 $D=1
M2342 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=202795 $Y=1334 $D=1
M2343 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=203275 $Y=-6292 $D=1
M2344 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=203485 $Y=1334 $D=1
M2345 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=203965 $Y=-6292 $D=1
M2346 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=204175 $Y=1334 $D=1
M2347 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=204655 $Y=-6292 $D=1
M2348 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=204865 $Y=1334 $D=1
M2349 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=205345 $Y=-6292 $D=1
M2350 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=205555 $Y=1334 $D=1
M2351 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=206035 $Y=-6292 $D=1
M2352 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=206245 $Y=1334 $D=1
M2353 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=206725 $Y=-6292 $D=1
M2354 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=206935 $Y=1334 $D=1
M2355 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=207415 $Y=-6292 $D=1
M2356 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=207625 $Y=1334 $D=1
M2357 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=208105 $Y=-6292 $D=1
M2358 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=208315 $Y=1334 $D=1
M2359 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=208795 $Y=-6292 $D=1
M2360 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=209005 $Y=1334 $D=1
M2361 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=209485 $Y=-6292 $D=1
M2362 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=209695 $Y=1334 $D=1
M2363 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=210175 $Y=-6292 $D=1
M2364 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=210385 $Y=1334 $D=1
M2365 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=210865 $Y=-6292 $D=1
M2366 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=211075 $Y=1334 $D=1
M2367 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=211555 $Y=-6292 $D=1
M2368 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=211765 $Y=1334 $D=1
M2369 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=212245 $Y=-6292 $D=1
M2370 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=212455 $Y=1334 $D=1
M2371 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=212935 $Y=-6292 $D=1
M2372 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=213145 $Y=1334 $D=1
M2373 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=213625 $Y=-6292 $D=1
M2374 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=213835 $Y=1334 $D=1
M2375 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=214315 $Y=-6292 $D=1
M2376 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=214525 $Y=1334 $D=1
M2377 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=215005 $Y=-6292 $D=1
M2378 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=215215 $Y=1334 $D=1
M2379 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=215695 $Y=-6292 $D=1
M2380 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=215905 $Y=1334 $D=1
M2381 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=216385 $Y=-6292 $D=1
M2382 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=216595 $Y=1334 $D=1
M2383 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=217075 $Y=-6292 $D=1
M2384 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=217285 $Y=1334 $D=1
M2385 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=217765 $Y=-6292 $D=1
M2386 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=217975 $Y=1334 $D=1
M2387 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=218455 $Y=-6292 $D=1
M2388 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=218665 $Y=1334 $D=1
M2389 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=219145 $Y=-6292 $D=1
M2390 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=219355 $Y=1334 $D=1
M2391 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=219835 $Y=-6292 $D=1
M2392 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=220045 $Y=1334 $D=1
M2393 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=220525 $Y=-6292 $D=1
M2394 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=220735 $Y=1334 $D=1
M2395 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=221215 $Y=-6292 $D=1
M2396 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=221425 $Y=1334 $D=1
M2397 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=221905 $Y=-6292 $D=1
M2398 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=222115 $Y=1334 $D=1
M2399 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=222595 $Y=-6292 $D=1
M2400 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=222805 $Y=1334 $D=1
M2401 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=223285 $Y=-6292 $D=1
M2402 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=223495 $Y=1334 $D=1
M2403 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=223975 $Y=-6292 $D=1
M2404 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=224185 $Y=1334 $D=1
M2405 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=224665 $Y=-6292 $D=1
M2406 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=224875 $Y=1334 $D=1
M2407 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=225355 $Y=-6292 $D=1
M2408 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=225565 $Y=1334 $D=1
M2409 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=226045 $Y=-6292 $D=1
M2410 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=226255 $Y=1334 $D=1
M2411 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=226735 $Y=-6292 $D=1
M2412 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=226945 $Y=1334 $D=1
M2413 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=227425 $Y=-6292 $D=1
M2414 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=227635 $Y=1334 $D=1
M2415 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=228115 $Y=-6292 $D=1
M2416 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=228325 $Y=1334 $D=1
M2417 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=228805 $Y=-6292 $D=1
M2418 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=229015 $Y=1334 $D=1
M2419 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=229495 $Y=-6292 $D=1
M2420 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=229705 $Y=1334 $D=1
M2421 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=230185 $Y=-6292 $D=1
M2422 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=230395 $Y=1334 $D=1
M2423 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=230875 $Y=-6292 $D=1
M2424 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=231085 $Y=1334 $D=1
M2425 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=231565 $Y=-6292 $D=1
M2426 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=231775 $Y=1334 $D=1
M2427 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=232255 $Y=-6292 $D=1
M2428 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=232465 $Y=1334 $D=1
M2429 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=232945 $Y=-6292 $D=1
M2430 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=233155 $Y=1334 $D=1
M2431 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=233635 $Y=-6292 $D=1
M2432 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=233845 $Y=1334 $D=1
M2433 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=234325 $Y=-6292 $D=1
M2434 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=234535 $Y=1334 $D=1
M2435 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=235015 $Y=-6292 $D=1
M2436 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=235225 $Y=1334 $D=1
M2437 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=235705 $Y=-6292 $D=1
M2438 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=235915 $Y=1334 $D=1
M2439 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=236395 $Y=-6292 $D=1
M2440 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=236605 $Y=1334 $D=1
M2441 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=237085 $Y=-6292 $D=1
M2442 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=237295 $Y=1334 $D=1
M2443 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=237775 $Y=-6292 $D=1
M2444 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=237985 $Y=1334 $D=1
M2445 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=238465 $Y=-6292 $D=1
M2446 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=238675 $Y=1334 $D=1
M2447 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=239155 $Y=-6292 $D=1
M2448 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=239365 $Y=1334 $D=1
M2449 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=5.2611e-13 AS=4.7073e-13 PD=5.7e-07 PS=5.1e-07 $X=239845 $Y=-6292 $D=1
M2450 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=240055 $Y=1334 $D=1
M2451 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=5.2611e-13 PD=5.1e-07 PS=5.7e-07 $X=240595 $Y=-6292 $D=1
M2452 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=240745 $Y=1334 $D=1
M2453 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=241285 $Y=-6292 $D=1
M2454 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=241435 $Y=1334 $D=1
M2455 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=241975 $Y=-6292 $D=1
M2456 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=242125 $Y=1334 $D=1
M2457 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=242665 $Y=-6292 $D=1
M2458 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=242815 $Y=1334 $D=1
M2459 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=243355 $Y=-6292 $D=1
M2460 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=243505 $Y=1334 $D=1
M2461 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=244045 $Y=-6292 $D=1
M2462 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=244195 $Y=1334 $D=1
M2463 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=244735 $Y=-6292 $D=1
M2464 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=244885 $Y=1334 $D=1
M2465 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=245425 $Y=-6292 $D=1
M2466 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=245575 $Y=1334 $D=1
M2467 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=246115 $Y=-6292 $D=1
M2468 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=246265 $Y=1334 $D=1
M2469 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=246805 $Y=-6292 $D=1
M2470 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=246955 $Y=1334 $D=1
M2471 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=247495 $Y=-6292 $D=1
M2472 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=247645 $Y=1334 $D=1
M2473 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=248185 $Y=-6292 $D=1
M2474 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=248335 $Y=1334 $D=1
M2475 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=248875 $Y=-6292 $D=1
M2476 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=249025 $Y=1334 $D=1
M2477 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=249565 $Y=-6292 $D=1
M2478 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=249715 $Y=1334 $D=1
M2479 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=250255 $Y=-6292 $D=1
M2480 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=250405 $Y=1334 $D=1
M2481 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=250945 $Y=-6292 $D=1
M2482 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=251095 $Y=1334 $D=1
M2483 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=251635 $Y=-6292 $D=1
M2484 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=251785 $Y=1334 $D=1
M2485 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=252325 $Y=-6292 $D=1
M2486 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=252475 $Y=1334 $D=1
M2487 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=253015 $Y=-6292 $D=1
M2488 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=253165 $Y=1334 $D=1
M2489 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=253705 $Y=-6292 $D=1
M2490 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=253855 $Y=1334 $D=1
M2491 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=254395 $Y=-6292 $D=1
M2492 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=254545 $Y=1334 $D=1
M2493 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=255085 $Y=-6292 $D=1
M2494 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=255235 $Y=1334 $D=1
M2495 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=255775 $Y=-6292 $D=1
M2496 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=255925 $Y=1334 $D=1
M2497 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=256465 $Y=-6292 $D=1
M2498 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=256615 $Y=1334 $D=1
M2499 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=257155 $Y=-6292 $D=1
M2500 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=257305 $Y=1334 $D=1
M2501 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=257845 $Y=-6292 $D=1
M2502 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=257995 $Y=1334 $D=1
M2503 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=258535 $Y=-6292 $D=1
M2504 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=258685 $Y=1334 $D=1
M2505 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=259225 $Y=-6292 $D=1
M2506 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=259375 $Y=1334 $D=1
M2507 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=259915 $Y=-6292 $D=1
M2508 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=260065 $Y=1334 $D=1
M2509 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=260605 $Y=-6292 $D=1
M2510 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=260755 $Y=1334 $D=1
M2511 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=261295 $Y=-6292 $D=1
M2512 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=261445 $Y=1334 $D=1
M2513 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=261985 $Y=-6292 $D=1
M2514 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=262135 $Y=1334 $D=1
M2515 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=262675 $Y=-6292 $D=1
M2516 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=262825 $Y=1334 $D=1
M2517 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=263365 $Y=-6292 $D=1
M2518 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=263515 $Y=1334 $D=1
M2519 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=264055 $Y=-6292 $D=1
M2520 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=264205 $Y=1334 $D=1
M2521 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=264745 $Y=-6292 $D=1
M2522 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=264895 $Y=1334 $D=1
M2523 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=265435 $Y=-6292 $D=1
M2524 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=265585 $Y=1334 $D=1
M2525 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=266125 $Y=-6292 $D=1
M2526 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=266275 $Y=1334 $D=1
M2527 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=266815 $Y=-6292 $D=1
M2528 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=266965 $Y=1334 $D=1
M2529 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=267505 $Y=-6292 $D=1
M2530 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=267655 $Y=1334 $D=1
M2531 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=268195 $Y=-6292 $D=1
M2532 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=268345 $Y=1334 $D=1
M2533 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=268885 $Y=-6292 $D=1
M2534 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=269035 $Y=1334 $D=1
M2535 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=269575 $Y=-6292 $D=1
M2536 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=269725 $Y=1334 $D=1
M2537 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=270265 $Y=-6292 $D=1
M2538 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=270415 $Y=1334 $D=1
M2539 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=270955 $Y=-6292 $D=1
M2540 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=271105 $Y=1334 $D=1
M2541 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=271645 $Y=-6292 $D=1
M2542 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=271795 $Y=1334 $D=1
M2543 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=272335 $Y=-6292 $D=1
M2544 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=272485 $Y=1334 $D=1
M2545 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=273025 $Y=-6292 $D=1
M2546 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=273175 $Y=1334 $D=1
M2547 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=273715 $Y=-6292 $D=1
M2548 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=273865 $Y=1334 $D=1
M2549 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=274405 $Y=-6292 $D=1
M2550 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=274555 $Y=1334 $D=1
M2551 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=275095 $Y=-6292 $D=1
M2552 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=275245 $Y=1334 $D=1
M2553 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=275785 $Y=-6292 $D=1
M2554 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=275935 $Y=1334 $D=1
M2555 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=276475 $Y=-6292 $D=1
M2556 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=276625 $Y=1334 $D=1
M2557 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=277165 $Y=-6292 $D=1
M2558 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=277315 $Y=1334 $D=1
M2559 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=277855 $Y=-6292 $D=1
M2560 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=278005 $Y=1334 $D=1
M2561 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=278545 $Y=-6292 $D=1
M2562 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=278695 $Y=1334 $D=1
M2563 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=279235 $Y=-6292 $D=1
M2564 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=279385 $Y=1334 $D=1
M2565 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=279925 $Y=-6292 $D=1
M2566 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=280075 $Y=1334 $D=1
M2567 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=280615 $Y=-6292 $D=1
M2568 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=280765 $Y=1334 $D=1
M2569 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=281305 $Y=-6292 $D=1
M2570 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=281455 $Y=1334 $D=1
M2571 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=281995 $Y=-6292 $D=1
M2572 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=282145 $Y=1334 $D=1
M2573 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=282685 $Y=-6292 $D=1
M2574 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=282835 $Y=1334 $D=1
M2575 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=283375 $Y=-6292 $D=1
M2576 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=283525 $Y=1334 $D=1
M2577 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=284065 $Y=-6292 $D=1
M2578 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=284215 $Y=1334 $D=1
M2579 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=284755 $Y=-6292 $D=1
M2580 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=284905 $Y=1334 $D=1
M2581 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=285445 $Y=-6292 $D=1
M2582 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=285595 $Y=1334 $D=1
M2583 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=286135 $Y=-6292 $D=1
M2584 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=286285 $Y=1334 $D=1
M2585 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=286825 $Y=-6292 $D=1
M2586 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=286975 $Y=1334 $D=1
M2587 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=287515 $Y=-6292 $D=1
M2588 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=287665 $Y=1334 $D=1
M2589 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=288205 $Y=-6292 $D=1
M2590 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=288355 $Y=1334 $D=1
M2591 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=288895 $Y=-6292 $D=1
M2592 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=289045 $Y=1334 $D=1
M2593 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=289585 $Y=-6292 $D=1
M2594 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=289735 $Y=1334 $D=1
M2595 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=290275 $Y=-6292 $D=1
M2596 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=290425 $Y=1334 $D=1
M2597 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=290965 $Y=-6292 $D=1
M2598 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=291115 $Y=1334 $D=1
M2599 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=291655 $Y=-6292 $D=1
M2600 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=291805 $Y=1334 $D=1
M2601 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=292345 $Y=-6292 $D=1
M2602 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=292495 $Y=1334 $D=1
M2603 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=293035 $Y=-6292 $D=1
M2604 VDD 15 Vbout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=293185 $Y=1334 $D=1
M2605 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=293725 $Y=-6292 $D=1
M2606 Vbout 15 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=293875 $Y=1334 $D=1
M2607 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=294415 $Y=-6292 $D=1
M2608 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=295105 $Y=-6292 $D=1
M2609 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=295795 $Y=-6292 $D=1
M2610 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=296485 $Y=-6292 $D=1
M2611 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=297175 $Y=-6292 $D=1
M2612 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=297865 $Y=-6292 $D=1
M2613 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=298555 $Y=-6292 $D=1
M2614 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=299245 $Y=-6292 $D=1
M2615 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=299935 $Y=-6292 $D=1
M2616 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=300625 $Y=-6292 $D=1
M2617 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=301315 $Y=-6292 $D=1
M2618 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=302005 $Y=-6292 $D=1
M2619 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=302695 $Y=-6292 $D=1
M2620 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=303385 $Y=-6292 $D=1
M2621 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=304075 $Y=-6292 $D=1
M2622 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=304765 $Y=-6292 $D=1
M2623 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=305455 $Y=-6292 $D=1
M2624 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=306145 $Y=-6292 $D=1
M2625 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=306835 $Y=-6292 $D=1
M2626 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=307525 $Y=-6292 $D=1
M2627 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=308215 $Y=-6292 $D=1
M2628 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=308905 $Y=-6292 $D=1
M2629 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=309595 $Y=-6292 $D=1
M2630 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=310285 $Y=-6292 $D=1
M2631 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=310975 $Y=-6292 $D=1
M2632 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=311665 $Y=-6292 $D=1
M2633 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=312355 $Y=-6292 $D=1
M2634 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=313045 $Y=-6292 $D=1
M2635 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=313735 $Y=-6292 $D=1
M2636 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=314425 $Y=-6292 $D=1
M2637 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=315115 $Y=-6292 $D=1
M2638 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=315805 $Y=-6292 $D=1
M2639 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=316495 $Y=-6292 $D=1
M2640 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=317185 $Y=-6292 $D=1
M2641 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=317875 $Y=-6292 $D=1
M2642 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=318565 $Y=-6292 $D=1
M2643 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=319255 $Y=-6292 $D=1
M2644 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=319945 $Y=-6292 $D=1
M2645 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=320635 $Y=-6292 $D=1
M2646 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=321325 $Y=-6292 $D=1
M2647 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=322015 $Y=-6292 $D=1
M2648 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=322705 $Y=-6292 $D=1
M2649 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=323395 $Y=-6292 $D=1
M2650 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=324085 $Y=-6292 $D=1
M2651 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=324775 $Y=-6292 $D=1
M2652 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=325465 $Y=-6292 $D=1
M2653 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=326155 $Y=-6292 $D=1
M2654 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=326845 $Y=-6292 $D=1
M2655 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=327535 $Y=-6292 $D=1
M2656 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=328225 $Y=-6292 $D=1
M2657 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=328915 $Y=-6292 $D=1
M2658 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=329605 $Y=-6292 $D=1
M2659 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=330295 $Y=-6292 $D=1
M2660 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=330985 $Y=-6292 $D=1
M2661 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=331675 $Y=-6292 $D=1
M2662 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=332365 $Y=-6292 $D=1
M2663 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=333055 $Y=-6292 $D=1
M2664 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=333745 $Y=-6292 $D=1
M2665 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=334435 $Y=-6292 $D=1
M2666 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=335125 $Y=-6292 $D=1
M2667 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=335815 $Y=-6292 $D=1
M2668 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=336505 $Y=-6292 $D=1
M2669 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=337195 $Y=-6292 $D=1
M2670 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=337885 $Y=-6292 $D=1
M2671 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=338575 $Y=-6292 $D=1
M2672 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=339265 $Y=-6292 $D=1
M2673 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=339955 $Y=-6292 $D=1
M2674 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=340645 $Y=-6292 $D=1
M2675 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=341335 $Y=-6292 $D=1
M2676 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=342025 $Y=-6292 $D=1
M2677 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=342715 $Y=-6292 $D=1
M2678 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=343405 $Y=-6292 $D=1
M2679 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=344095 $Y=-6292 $D=1
M2680 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=344785 $Y=-6292 $D=1
M2681 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=345475 $Y=-6292 $D=1
M2682 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=346165 $Y=-6292 $D=1
M2683 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=346855 $Y=-6292 $D=1
M2684 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=347545 $Y=-6292 $D=1
M2685 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=348235 $Y=-6292 $D=1
M2686 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=348925 $Y=-6292 $D=1
M2687 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=349615 $Y=-6292 $D=1
M2688 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=350305 $Y=-6292 $D=1
M2689 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=350995 $Y=-6292 $D=1
M2690 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=351685 $Y=-6292 $D=1
M2691 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=352375 $Y=-6292 $D=1
M2692 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=353065 $Y=-6292 $D=1
M2693 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=353755 $Y=-6292 $D=1
M2694 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=354445 $Y=-6292 $D=1
M2695 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=355135 $Y=-6292 $D=1
M2696 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=355825 $Y=-6292 $D=1
M2697 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=356515 $Y=-6292 $D=1
M2698 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=357205 $Y=-6292 $D=1
M2699 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=357895 $Y=-6292 $D=1
M2700 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=358585 $Y=-6292 $D=1
M2701 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=359275 $Y=-6292 $D=1
M2702 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=359965 $Y=-6292 $D=1
M2703 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=360655 $Y=-6292 $D=1
M2704 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=361345 $Y=-6292 $D=1
M2705 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=362035 $Y=-6292 $D=1
M2706 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=362725 $Y=-6292 $D=1
M2707 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=363415 $Y=-6292 $D=1
M2708 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=364105 $Y=-6292 $D=1
M2709 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=364795 $Y=-6292 $D=1
M2710 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=365485 $Y=-6292 $D=1
M2711 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=366175 $Y=-6292 $D=1
M2712 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=366865 $Y=-6292 $D=1
M2713 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=367555 $Y=-6292 $D=1
M2714 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=368245 $Y=-6292 $D=1
M2715 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=368935 $Y=-6292 $D=1
M2716 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=369625 $Y=-6292 $D=1
M2717 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=370315 $Y=-6292 $D=1
M2718 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=371005 $Y=-6292 $D=1
M2719 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=371695 $Y=-6292 $D=1
M2720 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=372385 $Y=-6292 $D=1
M2721 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=373075 $Y=-6292 $D=1
M2722 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=373765 $Y=-6292 $D=1
M2723 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=374455 $Y=-6292 $D=1
M2724 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=375145 $Y=-6292 $D=1
M2725 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=375835 $Y=-6292 $D=1
M2726 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=376525 $Y=-6292 $D=1
M2727 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=377215 $Y=-6292 $D=1
M2728 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=377905 $Y=-6292 $D=1
M2729 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=378595 $Y=-6292 $D=1
M2730 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=379285 $Y=-6292 $D=1
M2731 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=379975 $Y=-6292 $D=1
M2732 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=380665 $Y=-6292 $D=1
M2733 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=381355 $Y=-6292 $D=1
M2734 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=382045 $Y=-6292 $D=1
M2735 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=382735 $Y=-6292 $D=1
M2736 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=383425 $Y=-6292 $D=1
M2737 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=384115 $Y=-6292 $D=1
M2738 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=384805 $Y=-6292 $D=1
M2739 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=385495 $Y=-6292 $D=1
M2740 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=386185 $Y=-6292 $D=1
M2741 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=386875 $Y=-6292 $D=1
M2742 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=387565 $Y=-6292 $D=1
M2743 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=388255 $Y=-6292 $D=1
M2744 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=388945 $Y=-6292 $D=1
M2745 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=389635 $Y=-6292 $D=1
M2746 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=390325 $Y=-6292 $D=1
M2747 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=391015 $Y=-6292 $D=1
M2748 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=391705 $Y=-6292 $D=1
M2749 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=392395 $Y=-6292 $D=1
M2750 VDD 17 19 VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=393085 $Y=-6292 $D=1
M2751 19 17 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=393775 $Y=-6292 $D=1
M2752 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=9.0454e-13 PD=5.1e-07 PS=2.826e-06 $X=395335 $Y=-6292 $D=1
M2753 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=396025 $Y=-6292 $D=1
M2754 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=396715 $Y=-6292 $D=1
M2755 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=397405 $Y=-6292 $D=1
M2756 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=398095 $Y=-6292 $D=1
M2757 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=398785 $Y=-6292 $D=1
M2758 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=399475 $Y=-6292 $D=1
M2759 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=400165 $Y=-6292 $D=1
M2760 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=400855 $Y=-6292 $D=1
M2761 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=401545 $Y=-6292 $D=1
M2762 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=402235 $Y=-6292 $D=1
M2763 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=402925 $Y=-6292 $D=1
M2764 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=403615 $Y=-6292 $D=1
M2765 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=404305 $Y=-6292 $D=1
M2766 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=404995 $Y=-6292 $D=1
M2767 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=405685 $Y=-6292 $D=1
M2768 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=406375 $Y=-6292 $D=1
M2769 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=407065 $Y=-6292 $D=1
M2770 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=407755 $Y=-6292 $D=1
M2771 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=408445 $Y=-6292 $D=1
M2772 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=409135 $Y=-6292 $D=1
M2773 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=409825 $Y=-6292 $D=1
M2774 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=410515 $Y=-6292 $D=1
M2775 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=411205 $Y=-6292 $D=1
M2776 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=411895 $Y=-6292 $D=1
M2777 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=412585 $Y=-6292 $D=1
M2778 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=413275 $Y=-6292 $D=1
M2779 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=413965 $Y=-6292 $D=1
M2780 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=414655 $Y=-6292 $D=1
M2781 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=415345 $Y=-6292 $D=1
M2782 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=416035 $Y=-6292 $D=1
M2783 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=416725 $Y=-6292 $D=1
M2784 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=417415 $Y=-6292 $D=1
M2785 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=418105 $Y=-6292 $D=1
M2786 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=418795 $Y=-6292 $D=1
M2787 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=419485 $Y=-6292 $D=1
M2788 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=420175 $Y=-6292 $D=1
M2789 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=420865 $Y=-6292 $D=1
M2790 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=421555 $Y=-6292 $D=1
M2791 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=422245 $Y=-6292 $D=1
M2792 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=422935 $Y=-6292 $D=1
M2793 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=423625 $Y=-6292 $D=1
M2794 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=424315 $Y=-6292 $D=1
M2795 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=425005 $Y=-6292 $D=1
M2796 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=425695 $Y=-6292 $D=1
M2797 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=426385 $Y=-6292 $D=1
M2798 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=427075 $Y=-6292 $D=1
M2799 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=427765 $Y=-6292 $D=1
M2800 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=428455 $Y=-6292 $D=1
M2801 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=429145 $Y=-6292 $D=1
M2802 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=429835 $Y=-6292 $D=1
M2803 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=430525 $Y=-6292 $D=1
M2804 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=431215 $Y=-6292 $D=1
M2805 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=431905 $Y=-6292 $D=1
M2806 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=432595 $Y=-6292 $D=1
M2807 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=433285 $Y=-6292 $D=1
M2808 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=433975 $Y=-6292 $D=1
M2809 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=434665 $Y=-6292 $D=1
M2810 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=435355 $Y=-6292 $D=1
M2811 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=436045 $Y=-6292 $D=1
M2812 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=436735 $Y=-6292 $D=1
M2813 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=437425 $Y=-6292 $D=1
M2814 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=438115 $Y=-6292 $D=1
M2815 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=438805 $Y=-6292 $D=1
M2816 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=439495 $Y=-6292 $D=1
M2817 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=440185 $Y=-6292 $D=1
M2818 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=440875 $Y=-6292 $D=1
M2819 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=441565 $Y=-6292 $D=1
M2820 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=442255 $Y=-6292 $D=1
M2821 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=442945 $Y=-6292 $D=1
M2822 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=443635 $Y=-6292 $D=1
M2823 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=444325 $Y=-6292 $D=1
M2824 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=445015 $Y=-6292 $D=1
M2825 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=445705 $Y=-6292 $D=1
M2826 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=446395 $Y=-6292 $D=1
M2827 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=447085 $Y=-6292 $D=1
M2828 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=447775 $Y=-6292 $D=1
M2829 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=448465 $Y=-6292 $D=1
M2830 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=449155 $Y=-6292 $D=1
M2831 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=449845 $Y=-6292 $D=1
M2832 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=450535 $Y=-6292 $D=1
M2833 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=451225 $Y=-6292 $D=1
M2834 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=451915 $Y=-6292 $D=1
M2835 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=452605 $Y=-6292 $D=1
M2836 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=453295 $Y=-6292 $D=1
M2837 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=453985 $Y=-6292 $D=1
M2838 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=454675 $Y=-6292 $D=1
M2839 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=455365 $Y=-6292 $D=1
M2840 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=456055 $Y=-6292 $D=1
M2841 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=5.2611e-13 AS=4.7073e-13 PD=5.7e-07 PS=5.1e-07 $X=456745 $Y=-6292 $D=1
M2842 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=5.2611e-13 PD=5.1e-07 PS=5.7e-07 $X=457495 $Y=-6292 $D=1
M2843 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=458185 $Y=-6292 $D=1
M2844 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=458875 $Y=-6292 $D=1
M2845 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=459565 $Y=-6292 $D=1
M2846 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=460255 $Y=-6292 $D=1
M2847 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=460945 $Y=-6292 $D=1
M2848 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=461635 $Y=-6292 $D=1
M2849 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=462325 $Y=-6292 $D=1
M2850 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=463015 $Y=-6292 $D=1
M2851 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=463705 $Y=-6292 $D=1
M2852 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=464395 $Y=-6292 $D=1
M2853 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=465085 $Y=-6292 $D=1
M2854 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=465775 $Y=-6292 $D=1
M2855 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=466465 $Y=-6292 $D=1
M2856 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=467155 $Y=-6292 $D=1
M2857 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=467845 $Y=-6292 $D=1
M2858 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=468535 $Y=-6292 $D=1
M2859 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=469225 $Y=-6292 $D=1
M2860 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=469915 $Y=-6292 $D=1
M2861 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=470605 $Y=-6292 $D=1
M2862 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=471295 $Y=-6292 $D=1
M2863 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=471985 $Y=-6292 $D=1
M2864 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=472675 $Y=-6292 $D=1
M2865 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=473365 $Y=-6292 $D=1
M2866 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=474055 $Y=-6292 $D=1
M2867 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=474745 $Y=-6292 $D=1
M2868 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=475435 $Y=-6292 $D=1
M2869 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=476125 $Y=-6292 $D=1
M2870 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=476815 $Y=-6292 $D=1
M2871 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=477505 $Y=-6292 $D=1
M2872 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=478195 $Y=-6292 $D=1
M2873 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=478885 $Y=-6292 $D=1
M2874 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=479575 $Y=-6292 $D=1
M2875 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=480265 $Y=-6292 $D=1
M2876 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=480955 $Y=-6292 $D=1
M2877 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=481645 $Y=-6292 $D=1
M2878 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=482335 $Y=-6292 $D=1
M2879 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=483025 $Y=-6292 $D=1
M2880 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=483715 $Y=-6292 $D=1
M2881 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=484405 $Y=-6292 $D=1
M2882 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=485095 $Y=-6292 $D=1
M2883 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=485785 $Y=-6292 $D=1
M2884 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=486475 $Y=-6292 $D=1
M2885 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=487165 $Y=-6292 $D=1
M2886 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=487855 $Y=-6292 $D=1
M2887 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=488545 $Y=-6292 $D=1
M2888 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=489235 $Y=-6292 $D=1
M2889 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=489925 $Y=-6292 $D=1
M2890 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=490615 $Y=-6292 $D=1
M2891 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=491305 $Y=-6292 $D=1
M2892 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=491995 $Y=-6292 $D=1
M2893 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=492685 $Y=-6292 $D=1
M2894 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=493375 $Y=-6292 $D=1
M2895 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=494065 $Y=-6292 $D=1
M2896 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=494755 $Y=-6292 $D=1
M2897 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=495445 $Y=-6292 $D=1
M2898 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=496135 $Y=-6292 $D=1
M2899 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=496825 $Y=-6292 $D=1
M2900 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=497515 $Y=-6292 $D=1
M2901 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=498205 $Y=-6292 $D=1
M2902 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=498895 $Y=-6292 $D=1
M2903 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=499585 $Y=-6292 $D=1
M2904 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=500275 $Y=-6292 $D=1
M2905 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=500965 $Y=-6292 $D=1
M2906 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=501655 $Y=-6292 $D=1
M2907 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=502345 $Y=-6292 $D=1
M2908 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=503035 $Y=-6292 $D=1
M2909 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=503725 $Y=-6292 $D=1
M2910 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=504415 $Y=-6292 $D=1
M2911 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=505105 $Y=-6292 $D=1
M2912 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=505795 $Y=-6292 $D=1
M2913 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=506485 $Y=-6292 $D=1
M2914 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=507175 $Y=-6292 $D=1
M2915 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=507865 $Y=-6292 $D=1
M2916 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=508555 $Y=-6292 $D=1
M2917 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=509245 $Y=-6292 $D=1
M2918 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=509935 $Y=-6292 $D=1
M2919 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=510625 $Y=-6292 $D=1
M2920 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=511315 $Y=-6292 $D=1
M2921 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=512005 $Y=-6292 $D=1
M2922 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=512695 $Y=-6292 $D=1
M2923 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=513385 $Y=-6292 $D=1
M2924 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=514075 $Y=-6292 $D=1
M2925 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=514765 $Y=-6292 $D=1
M2926 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=515455 $Y=-6292 $D=1
M2927 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=516145 $Y=-6292 $D=1
M2928 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=516835 $Y=-6292 $D=1
M2929 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=517525 $Y=-6292 $D=1
M2930 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=518215 $Y=-6292 $D=1
M2931 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=518905 $Y=-6292 $D=1
M2932 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=519595 $Y=-6292 $D=1
M2933 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=520285 $Y=-6292 $D=1
M2934 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=520975 $Y=-6292 $D=1
M2935 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=521665 $Y=-6292 $D=1
M2936 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=522355 $Y=-6292 $D=1
M2937 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=523045 $Y=-6292 $D=1
M2938 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=523735 $Y=-6292 $D=1
M2939 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=524425 $Y=-6292 $D=1
M2940 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=525115 $Y=-6292 $D=1
M2941 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=525805 $Y=-6292 $D=1
M2942 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=526495 $Y=-6292 $D=1
M2943 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=527185 $Y=-6292 $D=1
M2944 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=527875 $Y=-6292 $D=1
M2945 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=528565 $Y=-6292 $D=1
M2946 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=529255 $Y=-6292 $D=1
M2947 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=529945 $Y=-6292 $D=1
M2948 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=530635 $Y=-6292 $D=1
M2949 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=531325 $Y=-6292 $D=1
M2950 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=532015 $Y=-6292 $D=1
M2951 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=532705 $Y=-6292 $D=1
M2952 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=533395 $Y=-6292 $D=1
M2953 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=534085 $Y=-6292 $D=1
M2954 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=534775 $Y=-6292 $D=1
M2955 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=535465 $Y=-6292 $D=1
M2956 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=536155 $Y=-6292 $D=1
M2957 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=536845 $Y=-6292 $D=1
M2958 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=537535 $Y=-6292 $D=1
M2959 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=538225 $Y=-6292 $D=1
M2960 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=538915 $Y=-6292 $D=1
M2961 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=539605 $Y=-6292 $D=1
M2962 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=540295 $Y=-6292 $D=1
M2963 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=540985 $Y=-6292 $D=1
M2964 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=541675 $Y=-6292 $D=1
M2965 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=542365 $Y=-6292 $D=1
M2966 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=543055 $Y=-6292 $D=1
M2967 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=543745 $Y=-6292 $D=1
M2968 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=544435 $Y=-6292 $D=1
M2969 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=545125 $Y=-6292 $D=1
M2970 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=545815 $Y=-6292 $D=1
M2971 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=546505 $Y=-6292 $D=1
M2972 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=547195 $Y=-6292 $D=1
M2973 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=547885 $Y=-6292 $D=1
M2974 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=548575 $Y=-6292 $D=1
M2975 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=549265 $Y=-6292 $D=1
M2976 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=549955 $Y=-6292 $D=1
M2977 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=550645 $Y=-6292 $D=1
M2978 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=551335 $Y=-6292 $D=1
M2979 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=552025 $Y=-6292 $D=1
M2980 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=552715 $Y=-6292 $D=1
M2981 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=553405 $Y=-6292 $D=1
M2982 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=554095 $Y=-6292 $D=1
M2983 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=554785 $Y=-6292 $D=1
M2984 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=555475 $Y=-6292 $D=1
M2985 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=556165 $Y=-6292 $D=1
M2986 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=556855 $Y=-6292 $D=1
M2987 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=557545 $Y=-6292 $D=1
M2988 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=558235 $Y=-6292 $D=1
M2989 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=558925 $Y=-6292 $D=1
M2990 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=559615 $Y=-6292 $D=1
M2991 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=560305 $Y=-6292 $D=1
M2992 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=560995 $Y=-6292 $D=1
M2993 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=561685 $Y=-6292 $D=1
M2994 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=562375 $Y=-6292 $D=1
M2995 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=563065 $Y=-6292 $D=1
M2996 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=563755 $Y=-6292 $D=1
M2997 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=564445 $Y=-6292 $D=1
M2998 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=565135 $Y=-6292 $D=1
M2999 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=565825 $Y=-6292 $D=1
M3000 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=566515 $Y=-6292 $D=1
M3001 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=567205 $Y=-6292 $D=1
M3002 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=567895 $Y=-6292 $D=1
M3003 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=568585 $Y=-6292 $D=1
M3004 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=569275 $Y=-6292 $D=1
M3005 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=569965 $Y=-6292 $D=1
M3006 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=570655 $Y=-6292 $D=1
M3007 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=571345 $Y=-6292 $D=1
M3008 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=572035 $Y=-6292 $D=1
M3009 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=572725 $Y=-6292 $D=1
M3010 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=573415 $Y=-6292 $D=1
M3011 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=574105 $Y=-6292 $D=1
M3012 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=574795 $Y=-6292 $D=1
M3013 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=575485 $Y=-6292 $D=1
M3014 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=576175 $Y=-6292 $D=1
M3015 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=576865 $Y=-6292 $D=1
M3016 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=577555 $Y=-6292 $D=1
M3017 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=578245 $Y=-6292 $D=1
M3018 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=578935 $Y=-6292 $D=1
M3019 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=579625 $Y=-6292 $D=1
M3020 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=580315 $Y=-6292 $D=1
M3021 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=581005 $Y=-6292 $D=1
M3022 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=581695 $Y=-6292 $D=1
M3023 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=582385 $Y=-6292 $D=1
M3024 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=583075 $Y=-6292 $D=1
M3025 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=583765 $Y=-6292 $D=1
M3026 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=584455 $Y=-6292 $D=1
M3027 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=585145 $Y=-6292 $D=1
M3028 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=585835 $Y=-6292 $D=1
M3029 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=586525 $Y=-6292 $D=1
M3030 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=587215 $Y=-6292 $D=1
M3031 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=587905 $Y=-6292 $D=1
M3032 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=588595 $Y=-6292 $D=1
M3033 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=589285 $Y=-6292 $D=1
M3034 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=589975 $Y=-6292 $D=1
M3035 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=590665 $Y=-6292 $D=1
M3036 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=591355 $Y=-6292 $D=1
M3037 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=592045 $Y=-6292 $D=1
M3038 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=592735 $Y=-6292 $D=1
M3039 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=593425 $Y=-6292 $D=1
M3040 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=594115 $Y=-6292 $D=1
M3041 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=594805 $Y=-6292 $D=1
M3042 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=595495 $Y=-6292 $D=1
M3043 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=596185 $Y=-6292 $D=1
M3044 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=596875 $Y=-6292 $D=1
M3045 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=597565 $Y=-6292 $D=1
M3046 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=598255 $Y=-6292 $D=1
M3047 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=598945 $Y=-6292 $D=1
M3048 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=599635 $Y=-6292 $D=1
M3049 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=600325 $Y=-6292 $D=1
M3050 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=601015 $Y=-6292 $D=1
M3051 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=601705 $Y=-6292 $D=1
M3052 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=602395 $Y=-6292 $D=1
M3053 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=603085 $Y=-6292 $D=1
M3054 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=603775 $Y=-6292 $D=1
M3055 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=604465 $Y=-6292 $D=1
M3056 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=605155 $Y=-6292 $D=1
M3057 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=605845 $Y=-6292 $D=1
M3058 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=606535 $Y=-6292 $D=1
M3059 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=607225 $Y=-6292 $D=1
M3060 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=607915 $Y=-6292 $D=1
M3061 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=608605 $Y=-6292 $D=1
M3062 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=609295 $Y=-6292 $D=1
M3063 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=609985 $Y=-6292 $D=1
M3064 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=610675 $Y=-6292 $D=1
M3065 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=611365 $Y=-6292 $D=1
M3066 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=612055 $Y=-6292 $D=1
M3067 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=612745 $Y=-6292 $D=1
M3068 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=613435 $Y=-6292 $D=1
M3069 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=614125 $Y=-6292 $D=1
M3070 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=614815 $Y=-6292 $D=1
M3071 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=615505 $Y=-6292 $D=1
M3072 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=616195 $Y=-6292 $D=1
M3073 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=616885 $Y=-6292 $D=1
M3074 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=617575 $Y=-6292 $D=1
M3075 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=618265 $Y=-6292 $D=1
M3076 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=618955 $Y=-6292 $D=1
M3077 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=619645 $Y=-6292 $D=1
M3078 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=620335 $Y=-6292 $D=1
M3079 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=621025 $Y=-6292 $D=1
M3080 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=621715 $Y=-6292 $D=1
M3081 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=622405 $Y=-6292 $D=1
M3082 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=623095 $Y=-6292 $D=1
M3083 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=623785 $Y=-6292 $D=1
M3084 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=624475 $Y=-6292 $D=1
M3085 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=625165 $Y=-6292 $D=1
M3086 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=625855 $Y=-6292 $D=1
M3087 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=626545 $Y=-6292 $D=1
M3088 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=627235 $Y=-6292 $D=1
M3089 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=627925 $Y=-6292 $D=1
M3090 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=628615 $Y=-6292 $D=1
M3091 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=629305 $Y=-6292 $D=1
M3092 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=629995 $Y=-6292 $D=1
M3093 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=630685 $Y=-6292 $D=1
M3094 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=631375 $Y=-6292 $D=1
M3095 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=632065 $Y=-6292 $D=1
M3096 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=632755 $Y=-6292 $D=1
M3097 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=633445 $Y=-6292 $D=1
M3098 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=634135 $Y=-6292 $D=1
M3099 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=634825 $Y=-6292 $D=1
M3100 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=635515 $Y=-6292 $D=1
M3101 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=636205 $Y=-6292 $D=1
M3102 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=636895 $Y=-6292 $D=1
M3103 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=637585 $Y=-6292 $D=1
M3104 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=638275 $Y=-6292 $D=1
M3105 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=638965 $Y=-6292 $D=1
M3106 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=639655 $Y=-6292 $D=1
M3107 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=640345 $Y=-6292 $D=1
M3108 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=641035 $Y=-6292 $D=1
M3109 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=641725 $Y=-6292 $D=1
M3110 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=642415 $Y=-6292 $D=1
M3111 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=643105 $Y=-6292 $D=1
M3112 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=643795 $Y=-6292 $D=1
M3113 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=644485 $Y=-6292 $D=1
M3114 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=645175 $Y=-6292 $D=1
M3115 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=645865 $Y=-6292 $D=1
M3116 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=646555 $Y=-6292 $D=1
M3117 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=647245 $Y=-6292 $D=1
M3118 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=647935 $Y=-6292 $D=1
M3119 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=648625 $Y=-6292 $D=1
M3120 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=649315 $Y=-6292 $D=1
M3121 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=650005 $Y=-6292 $D=1
M3122 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=650695 $Y=-6292 $D=1
M3123 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=651385 $Y=-6292 $D=1
M3124 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=652075 $Y=-6292 $D=1
M3125 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=652765 $Y=-6292 $D=1
M3126 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=653455 $Y=-6292 $D=1
M3127 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=654145 $Y=-6292 $D=1
M3128 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=654835 $Y=-6292 $D=1
M3129 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=655525 $Y=-6292 $D=1
M3130 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=656215 $Y=-6292 $D=1
M3131 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=656905 $Y=-6292 $D=1
M3132 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=657595 $Y=-6292 $D=1
M3133 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=658285 $Y=-6292 $D=1
M3134 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=658975 $Y=-6292 $D=1
M3135 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=659665 $Y=-6292 $D=1
M3136 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=660355 $Y=-6292 $D=1
M3137 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=661045 $Y=-6292 $D=1
M3138 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=661735 $Y=-6292 $D=1
M3139 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=662425 $Y=-6292 $D=1
M3140 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=663115 $Y=-6292 $D=1
M3141 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=663805 $Y=-6292 $D=1
M3142 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=664495 $Y=-6292 $D=1
M3143 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=665185 $Y=-6292 $D=1
M3144 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=665875 $Y=-6292 $D=1
M3145 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=666565 $Y=-6292 $D=1
M3146 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=667255 $Y=-6292 $D=1
M3147 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=667945 $Y=-6292 $D=1
M3148 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=668635 $Y=-6292 $D=1
M3149 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=669325 $Y=-6292 $D=1
M3150 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=670015 $Y=-6292 $D=1
M3151 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=670705 $Y=-6292 $D=1
M3152 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=671395 $Y=-6292 $D=1
M3153 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=5.2611e-13 AS=4.7073e-13 PD=5.7e-07 PS=5.1e-07 $X=672085 $Y=-6292 $D=1
M3154 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=5.2611e-13 PD=5.1e-07 PS=5.7e-07 $X=672835 $Y=-6292 $D=1
M3155 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=673525 $Y=-6292 $D=1
M3156 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=674215 $Y=-6292 $D=1
M3157 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=674905 $Y=-6292 $D=1
M3158 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=675595 $Y=-6292 $D=1
M3159 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=676285 $Y=-6292 $D=1
M3160 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=676975 $Y=-6292 $D=1
M3161 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=677665 $Y=-6292 $D=1
M3162 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=678355 $Y=-6292 $D=1
M3163 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=679045 $Y=-6292 $D=1
M3164 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=679735 $Y=-6292 $D=1
M3165 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=680425 $Y=-6292 $D=1
M3166 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=681115 $Y=-6292 $D=1
M3167 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=681805 $Y=-6292 $D=1
M3168 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=682495 $Y=-6292 $D=1
M3169 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=683185 $Y=-6292 $D=1
M3170 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=683875 $Y=-6292 $D=1
M3171 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=684565 $Y=-6292 $D=1
M3172 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=685255 $Y=-6292 $D=1
M3173 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=685945 $Y=-6292 $D=1
M3174 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=686635 $Y=-6292 $D=1
M3175 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=687325 $Y=-6292 $D=1
M3176 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=688015 $Y=-6292 $D=1
M3177 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=688705 $Y=-6292 $D=1
M3178 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=689395 $Y=-6292 $D=1
M3179 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=690085 $Y=-6292 $D=1
M3180 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=690775 $Y=-6292 $D=1
M3181 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=691465 $Y=-6292 $D=1
M3182 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=692155 $Y=-6292 $D=1
M3183 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=692845 $Y=-6292 $D=1
M3184 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=693535 $Y=-6292 $D=1
M3185 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=694225 $Y=-6292 $D=1
M3186 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=694915 $Y=-6292 $D=1
M3187 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=695605 $Y=-6292 $D=1
M3188 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=696295 $Y=-6292 $D=1
M3189 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=696985 $Y=-6292 $D=1
M3190 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=697675 $Y=-6292 $D=1
M3191 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=698365 $Y=-6292 $D=1
M3192 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=699055 $Y=-6292 $D=1
M3193 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=699745 $Y=-6292 $D=1
M3194 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=700435 $Y=-6292 $D=1
M3195 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=701125 $Y=-6292 $D=1
M3196 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=701815 $Y=-6292 $D=1
M3197 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=702505 $Y=-6292 $D=1
M3198 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=703195 $Y=-6292 $D=1
M3199 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=703885 $Y=-6292 $D=1
M3200 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=704575 $Y=-6292 $D=1
M3201 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=705265 $Y=-6292 $D=1
M3202 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=705955 $Y=-6292 $D=1
M3203 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=706645 $Y=-6292 $D=1
M3204 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=707335 $Y=-6292 $D=1
M3205 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=708025 $Y=-6292 $D=1
M3206 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=708715 $Y=-6292 $D=1
M3207 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=709405 $Y=-6292 $D=1
M3208 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=710095 $Y=-6292 $D=1
M3209 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=710785 $Y=-6292 $D=1
M3210 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=711475 $Y=-6292 $D=1
M3211 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=712165 $Y=-6292 $D=1
M3212 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=712855 $Y=-6292 $D=1
M3213 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=713545 $Y=-6292 $D=1
M3214 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=714235 $Y=-6292 $D=1
M3215 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=714925 $Y=-6292 $D=1
M3216 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=715615 $Y=-6292 $D=1
M3217 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=716305 $Y=-6292 $D=1
M3218 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=716995 $Y=-6292 $D=1
M3219 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=717685 $Y=-6292 $D=1
M3220 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=718375 $Y=-6292 $D=1
M3221 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=719065 $Y=-6292 $D=1
M3222 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=719755 $Y=-6292 $D=1
M3223 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=720445 $Y=-6292 $D=1
M3224 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=721135 $Y=-6292 $D=1
M3225 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=721825 $Y=-6292 $D=1
M3226 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=722515 $Y=-6292 $D=1
M3227 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=723205 $Y=-6292 $D=1
M3228 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=723895 $Y=-6292 $D=1
M3229 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=724585 $Y=-6292 $D=1
M3230 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=725275 $Y=-6292 $D=1
M3231 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=725965 $Y=-6292 $D=1
M3232 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=726655 $Y=-6292 $D=1
M3233 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=727345 $Y=-6292 $D=1
M3234 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=728035 $Y=-6292 $D=1
M3235 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=728725 $Y=-6292 $D=1
M3236 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=729415 $Y=-6292 $D=1
M3237 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=730105 $Y=-6292 $D=1
M3238 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=730795 $Y=-6292 $D=1
M3239 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=731485 $Y=-6292 $D=1
M3240 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=732175 $Y=-6292 $D=1
M3241 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=732865 $Y=-6292 $D=1
M3242 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=733555 $Y=-6292 $D=1
M3243 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=734245 $Y=-6292 $D=1
M3244 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=734935 $Y=-6292 $D=1
M3245 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=735625 $Y=-6292 $D=1
M3246 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=736315 $Y=-6292 $D=1
M3247 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=737005 $Y=-6292 $D=1
M3248 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=737695 $Y=-6292 $D=1
M3249 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=738385 $Y=-6292 $D=1
M3250 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=739075 $Y=-6292 $D=1
M3251 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=739765 $Y=-6292 $D=1
M3252 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=740455 $Y=-6292 $D=1
M3253 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=741145 $Y=-6292 $D=1
M3254 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=741835 $Y=-6292 $D=1
M3255 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=742525 $Y=-6292 $D=1
M3256 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=743215 $Y=-6292 $D=1
M3257 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=743905 $Y=-6292 $D=1
M3258 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=744595 $Y=-6292 $D=1
M3259 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=745285 $Y=-6292 $D=1
M3260 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=745975 $Y=-6292 $D=1
M3261 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=746665 $Y=-6292 $D=1
M3262 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=747355 $Y=-6292 $D=1
M3263 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=748045 $Y=-6292 $D=1
M3264 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=748735 $Y=-6292 $D=1
M3265 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=749425 $Y=-6292 $D=1
M3266 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=750115 $Y=-6292 $D=1
M3267 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=750805 $Y=-6292 $D=1
M3268 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=751495 $Y=-6292 $D=1
M3269 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=752185 $Y=-6292 $D=1
M3270 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=752875 $Y=-6292 $D=1
M3271 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=753565 $Y=-6292 $D=1
M3272 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=754255 $Y=-6292 $D=1
M3273 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=754945 $Y=-6292 $D=1
M3274 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=755635 $Y=-6292 $D=1
M3275 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=756325 $Y=-6292 $D=1
M3276 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=757015 $Y=-6292 $D=1
M3277 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=757705 $Y=-6292 $D=1
M3278 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=758395 $Y=-6292 $D=1
M3279 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=759085 $Y=-6292 $D=1
M3280 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=759775 $Y=-6292 $D=1
M3281 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=760465 $Y=-6292 $D=1
M3282 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=761155 $Y=-6292 $D=1
M3283 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=761845 $Y=-6292 $D=1
M3284 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=762535 $Y=-6292 $D=1
M3285 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=763225 $Y=-6292 $D=1
M3286 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=763915 $Y=-6292 $D=1
M3287 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=764605 $Y=-6292 $D=1
M3288 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=765295 $Y=-6292 $D=1
M3289 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=765985 $Y=-6292 $D=1
M3290 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=766675 $Y=-6292 $D=1
M3291 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=767365 $Y=-6292 $D=1
M3292 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=768055 $Y=-6292 $D=1
M3293 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=768745 $Y=-6292 $D=1
M3294 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=769435 $Y=-6292 $D=1
M3295 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=770125 $Y=-6292 $D=1
M3296 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=770815 $Y=-6292 $D=1
M3297 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=771505 $Y=-6292 $D=1
M3298 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=772195 $Y=-6292 $D=1
M3299 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=772885 $Y=-6292 $D=1
M3300 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=773575 $Y=-6292 $D=1
M3301 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=774265 $Y=-6292 $D=1
M3302 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=774955 $Y=-6292 $D=1
M3303 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=775645 $Y=-6292 $D=1
M3304 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=776335 $Y=-6292 $D=1
M3305 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=777025 $Y=-6292 $D=1
M3306 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=777715 $Y=-6292 $D=1
M3307 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=778405 $Y=-6292 $D=1
M3308 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=779095 $Y=-6292 $D=1
M3309 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=779785 $Y=-6292 $D=1
M3310 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=780475 $Y=-6292 $D=1
M3311 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=781165 $Y=-6292 $D=1
M3312 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=781855 $Y=-6292 $D=1
M3313 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=782545 $Y=-6292 $D=1
M3314 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=783235 $Y=-6292 $D=1
M3315 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=783925 $Y=-6292 $D=1
M3316 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=784615 $Y=-6292 $D=1
M3317 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=785305 $Y=-6292 $D=1
M3318 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=785995 $Y=-6292 $D=1
M3319 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=786685 $Y=-6292 $D=1
M3320 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=787375 $Y=-6292 $D=1
M3321 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=788065 $Y=-6292 $D=1
M3322 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=788755 $Y=-6292 $D=1
M3323 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=789445 $Y=-6292 $D=1
M3324 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=790135 $Y=-6292 $D=1
M3325 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=790825 $Y=-6292 $D=1
M3326 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=791515 $Y=-6292 $D=1
M3327 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=792205 $Y=-6292 $D=1
M3328 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=792895 $Y=-6292 $D=1
M3329 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=793585 $Y=-6292 $D=1
M3330 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=794275 $Y=-6292 $D=1
M3331 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=794965 $Y=-6292 $D=1
M3332 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=795655 $Y=-6292 $D=1
M3333 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=796345 $Y=-6292 $D=1
M3334 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=797035 $Y=-6292 $D=1
M3335 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=797725 $Y=-6292 $D=1
M3336 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=798415 $Y=-6292 $D=1
M3337 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=799105 $Y=-6292 $D=1
M3338 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=799795 $Y=-6292 $D=1
M3339 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=800485 $Y=-6292 $D=1
M3340 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=801175 $Y=-6292 $D=1
M3341 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=801865 $Y=-6292 $D=1
M3342 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=802555 $Y=-6292 $D=1
M3343 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=803245 $Y=-6292 $D=1
M3344 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=803935 $Y=-6292 $D=1
M3345 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=804625 $Y=-6292 $D=1
M3346 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=805315 $Y=-6292 $D=1
M3347 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=806005 $Y=-6292 $D=1
M3348 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=806695 $Y=-6292 $D=1
M3349 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=807385 $Y=-6292 $D=1
M3350 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=808075 $Y=-6292 $D=1
M3351 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=808765 $Y=-6292 $D=1
M3352 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=809455 $Y=-6292 $D=1
M3353 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=810145 $Y=-6292 $D=1
M3354 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=810835 $Y=-6292 $D=1
M3355 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=811525 $Y=-6292 $D=1
M3356 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=812215 $Y=-6292 $D=1
M3357 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=812905 $Y=-6292 $D=1
M3358 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=813595 $Y=-6292 $D=1
M3359 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=814285 $Y=-6292 $D=1
M3360 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=814975 $Y=-6292 $D=1
M3361 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=815665 $Y=-6292 $D=1
M3362 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=816355 $Y=-6292 $D=1
M3363 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=817045 $Y=-6292 $D=1
M3364 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=817735 $Y=-6292 $D=1
M3365 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=818425 $Y=-6292 $D=1
M3366 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=819115 $Y=-6292 $D=1
M3367 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=819805 $Y=-6292 $D=1
M3368 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=820495 $Y=-6292 $D=1
M3369 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=821185 $Y=-6292 $D=1
M3370 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=821875 $Y=-6292 $D=1
M3371 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=822565 $Y=-6292 $D=1
M3372 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=823255 $Y=-6292 $D=1
M3373 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=823945 $Y=-6292 $D=1
M3374 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=824635 $Y=-6292 $D=1
M3375 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=825325 $Y=-6292 $D=1
M3376 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=826015 $Y=-6292 $D=1
M3377 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=826705 $Y=-6292 $D=1
M3378 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=827395 $Y=-6292 $D=1
M3379 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=828085 $Y=-6292 $D=1
M3380 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=828775 $Y=-6292 $D=1
M3381 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=829465 $Y=-6292 $D=1
M3382 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=830155 $Y=-6292 $D=1
M3383 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=830845 $Y=-6292 $D=1
M3384 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=831535 $Y=-6292 $D=1
M3385 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=832225 $Y=-6292 $D=1
M3386 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=832915 $Y=-6292 $D=1
M3387 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=833605 $Y=-6292 $D=1
M3388 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=834295 $Y=-6292 $D=1
M3389 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=834985 $Y=-6292 $D=1
M3390 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=835675 $Y=-6292 $D=1
M3391 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=836365 $Y=-6292 $D=1
M3392 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=837055 $Y=-6292 $D=1
M3393 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=837745 $Y=-6292 $D=1
M3394 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=838435 $Y=-6292 $D=1
M3395 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=839125 $Y=-6292 $D=1
M3396 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=839815 $Y=-6292 $D=1
M3397 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=840505 $Y=-6292 $D=1
M3398 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=841195 $Y=-6292 $D=1
M3399 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=841885 $Y=-6292 $D=1
M3400 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=842575 $Y=-6292 $D=1
M3401 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=843265 $Y=-6292 $D=1
M3402 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=843955 $Y=-6292 $D=1
M3403 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=844645 $Y=-6292 $D=1
M3404 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=845335 $Y=-6292 $D=1
M3405 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=846025 $Y=-6292 $D=1
M3406 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=846715 $Y=-6292 $D=1
M3407 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=847405 $Y=-6292 $D=1
M3408 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=848095 $Y=-6292 $D=1
M3409 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=848785 $Y=-6292 $D=1
M3410 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=849475 $Y=-6292 $D=1
M3411 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=850165 $Y=-6292 $D=1
M3412 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=850855 $Y=-6292 $D=1
M3413 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=851545 $Y=-6292 $D=1
M3414 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=852235 $Y=-6292 $D=1
M3415 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=852925 $Y=-6292 $D=1
M3416 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=853615 $Y=-6292 $D=1
M3417 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=854305 $Y=-6292 $D=1
M3418 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=854995 $Y=-6292 $D=1
M3419 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=855685 $Y=-6292 $D=1
M3420 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=856375 $Y=-6292 $D=1
M3421 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=857065 $Y=-6292 $D=1
M3422 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=857755 $Y=-6292 $D=1
M3423 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=858445 $Y=-6292 $D=1
M3424 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=859135 $Y=-6292 $D=1
M3425 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=859825 $Y=-6292 $D=1
M3426 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=860515 $Y=-6292 $D=1
M3427 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=861205 $Y=-6292 $D=1
M3428 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=861895 $Y=-6292 $D=1
M3429 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=862585 $Y=-6292 $D=1
M3430 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=863275 $Y=-6292 $D=1
M3431 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=863965 $Y=-6292 $D=1
M3432 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=864655 $Y=-6292 $D=1
M3433 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=865345 $Y=-6292 $D=1
M3434 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=866035 $Y=-6292 $D=1
M3435 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=866725 $Y=-6292 $D=1
M3436 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=867415 $Y=-6292 $D=1
M3437 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=868105 $Y=-6292 $D=1
M3438 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=868795 $Y=-6292 $D=1
M3439 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=869485 $Y=-6292 $D=1
M3440 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=870175 $Y=-6292 $D=1
M3441 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=870865 $Y=-6292 $D=1
M3442 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=871555 $Y=-6292 $D=1
M3443 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=872245 $Y=-6292 $D=1
M3444 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=872935 $Y=-6292 $D=1
M3445 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=873625 $Y=-6292 $D=1
M3446 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=874315 $Y=-6292 $D=1
M3447 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=875005 $Y=-6292 $D=1
M3448 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=875695 $Y=-6292 $D=1
M3449 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=876385 $Y=-6292 $D=1
M3450 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=877075 $Y=-6292 $D=1
M3451 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=877765 $Y=-6292 $D=1
M3452 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=878455 $Y=-6292 $D=1
M3453 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=879145 $Y=-6292 $D=1
M3454 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=879835 $Y=-6292 $D=1
M3455 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=880525 $Y=-6292 $D=1
M3456 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=881215 $Y=-6292 $D=1
M3457 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=881905 $Y=-6292 $D=1
M3458 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=882595 $Y=-6292 $D=1
M3459 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=883285 $Y=-6292 $D=1
M3460 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=883975 $Y=-6292 $D=1
M3461 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=884665 $Y=-6292 $D=1
M3462 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=885355 $Y=-6292 $D=1
M3463 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=886045 $Y=-6292 $D=1
M3464 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=886735 $Y=-6292 $D=1
M3465 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=887425 $Y=-6292 $D=1
M3466 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=888115 $Y=-6292 $D=1
M3467 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=888805 $Y=-6292 $D=1
M3468 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=889495 $Y=-6292 $D=1
M3469 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=890185 $Y=-6292 $D=1
M3470 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=890875 $Y=-6292 $D=1
M3471 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=891565 $Y=-6292 $D=1
M3472 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=892255 $Y=-6292 $D=1
M3473 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=892945 $Y=-6292 $D=1
M3474 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=893635 $Y=-6292 $D=1
M3475 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=894325 $Y=-6292 $D=1
M3476 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=895015 $Y=-6292 $D=1
M3477 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=895705 $Y=-6292 $D=1
M3478 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=896395 $Y=-6292 $D=1
M3479 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=897085 $Y=-6292 $D=1
M3480 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=897775 $Y=-6292 $D=1
M3481 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=898465 $Y=-6292 $D=1
M3482 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=899155 $Y=-6292 $D=1
M3483 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=899845 $Y=-6292 $D=1
M3484 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=900535 $Y=-6292 $D=1
M3485 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=901225 $Y=-6292 $D=1
M3486 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=901915 $Y=-6292 $D=1
M3487 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=902605 $Y=-6292 $D=1
M3488 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=903295 $Y=-6292 $D=1
M3489 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=903985 $Y=-6292 $D=1
M3490 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=904675 $Y=-6292 $D=1
M3491 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=905365 $Y=-6292 $D=1
M3492 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=906055 $Y=-6292 $D=1
M3493 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=906745 $Y=-6292 $D=1
M3494 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=907435 $Y=-6292 $D=1
M3495 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=908125 $Y=-6292 $D=1
M3496 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=908815 $Y=-6292 $D=1
M3497 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=909505 $Y=-6292 $D=1
M3498 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=910195 $Y=-6292 $D=1
M3499 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=910885 $Y=-6292 $D=1
M3500 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=911575 $Y=-6292 $D=1
M3501 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=912265 $Y=-6292 $D=1
M3502 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=912955 $Y=-6292 $D=1
M3503 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=913645 $Y=-6292 $D=1
M3504 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=914335 $Y=-6292 $D=1
M3505 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=915025 $Y=-6292 $D=1
M3506 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=915715 $Y=-6292 $D=1
M3507 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=916405 $Y=-6292 $D=1
M3508 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=917095 $Y=-6292 $D=1
M3509 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=917785 $Y=-6292 $D=1
M3510 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=918475 $Y=-6292 $D=1
M3511 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=919165 $Y=-6292 $D=1
M3512 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=919855 $Y=-6292 $D=1
M3513 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=920545 $Y=-6292 $D=1
M3514 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=921235 $Y=-6292 $D=1
M3515 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=921925 $Y=-6292 $D=1
M3516 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=922615 $Y=-6292 $D=1
M3517 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=923305 $Y=-6292 $D=1
M3518 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=923995 $Y=-6292 $D=1
M3519 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=924685 $Y=-6292 $D=1
M3520 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=925375 $Y=-6292 $D=1
M3521 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=926065 $Y=-6292 $D=1
M3522 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=926755 $Y=-6292 $D=1
M3523 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=927445 $Y=-6292 $D=1
M3524 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=928135 $Y=-6292 $D=1
M3525 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=928825 $Y=-6292 $D=1
M3526 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=929515 $Y=-6292 $D=1
M3527 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=930205 $Y=-6292 $D=1
M3528 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=930895 $Y=-6292 $D=1
M3529 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=931585 $Y=-6292 $D=1
M3530 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=932275 $Y=-6292 $D=1
M3531 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=932965 $Y=-6292 $D=1
M3532 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=933655 $Y=-6292 $D=1
M3533 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=934345 $Y=-6292 $D=1
M3534 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=935035 $Y=-6292 $D=1
M3535 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=935725 $Y=-6292 $D=1
M3536 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=936415 $Y=-6292 $D=1
M3537 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=937105 $Y=-6292 $D=1
M3538 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=937795 $Y=-6292 $D=1
M3539 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=938485 $Y=-6292 $D=1
M3540 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=939175 $Y=-6292 $D=1
M3541 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=939865 $Y=-6292 $D=1
M3542 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=940555 $Y=-6292 $D=1
M3543 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=941245 $Y=-6292 $D=1
M3544 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=941935 $Y=-6292 $D=1
M3545 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=942625 $Y=-6292 $D=1
M3546 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=943315 $Y=-6292 $D=1
M3547 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=944005 $Y=-6292 $D=1
M3548 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=944695 $Y=-6292 $D=1
M3549 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=945385 $Y=-6292 $D=1
M3550 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=946075 $Y=-6292 $D=1
M3551 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=946765 $Y=-6292 $D=1
M3552 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=947455 $Y=-6292 $D=1
M3553 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=948145 $Y=-6292 $D=1
M3554 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=948835 $Y=-6292 $D=1
M3555 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=949525 $Y=-6292 $D=1
M3556 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=950215 $Y=-6292 $D=1
M3557 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=950905 $Y=-6292 $D=1
M3558 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=951595 $Y=-6292 $D=1
M3559 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=952285 $Y=-6292 $D=1
M3560 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=952975 $Y=-6292 $D=1
M3561 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=953665 $Y=-6292 $D=1
M3562 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=954355 $Y=-6292 $D=1
M3563 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=955045 $Y=-6292 $D=1
M3564 Vcout 19 VDD VDD P_18 L=1.8e-07 W=1.85e-06 AD=4.7073e-13 AS=4.7073e-13 PD=5.1e-07 PS=5.1e-07 $X=955735 $Y=-6292 $D=1
M3565 VDD 19 Vcout VDD P_18 L=1.8e-07 W=1.85e-06 AD=9.0454e-13 AS=4.7073e-13 PD=2.826e-06 PS=5.1e-07 $X=956425 $Y=-6292 $D=1
.ENDS
***************************************
