************************************************************************
* auCdl Netlist:
* 
* Library Name:  HW3
* Top Cell Name: SRL
* View Name:     schematic
* Netlisted on:  Nov 27 23:13:19 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: HW3
* Cell Name:    SRL
* View Name:    schematic
************************************************************************

.SUBCKT SRL CLK Q QB R S VDD VSS
*.PININFO R:I S:I Q:O QB:O CLK:B VDD:B VSS:B
MM5 Q QB VDD VDD p_18 W=500.00n L=180.00n m=1
MM4 QB Q VDD VDD p_18 W=500.00n L=180.00n m=1
MM3 Q QB VSS VSS n_18 W=500.0n L=180.00n m=1
MM2 QB Q VSS VSS n_18 W=500.0n L=180.00n m=1
MM1 S CLK Q VSS n_18 W=3.38U L=180.00n m=1
MM0 QB CLK R VSS n_18 W=3.38U L=180.00n m=1
.ENDS

